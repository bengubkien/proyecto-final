XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C��V->�/�n��� �#�� �w�H��m����tkz>����ƣ��%'#B���ͽVMIwԸ!}n��I��`bN�����k������S�,ӔU��$q�	���5����z�m3���J#͠f���T��,�<������4җEt�C)c*��Ђ��tDQx�fԄ�pkG$Î����D	wi��n�6�sa�����}��$�dj���Dɒ�a�w	���L�����nt@2)�dؠ�"�5b���ii:.��L����kU��Db_N���-y����֏[�cĉIӱ����2PGF���-�b U����:
��M�tH)��?�c�TQ-�g�Α.���'���P�̣�c��&�Q�)�n�	x�ٵ���>�����)DJ�H���pRj���a�"M�#͹�1<�q~l�%�?7�O��,��+���y|�h��p�C٪L�n�qvF4��3n����}��,	5���<�-W��C����/�le���;s}���ͧ��͸���=K�_*���~	S��'>�oeQƆe-����;����϶��WT� �L�`���D�}�~�j�Ts$|;����-i,T�,\'okG<U��]����϶�����f��[���=�*��u����q�t��#�=�w9e�<i)ab�Zk$(7���ck a�)s��G�M5��sk"r����W;�ۜ���.���r�a�0���.*�o�J �&}����9����W7u�,��,�Gm�{�X;��1=���~XlxVHYEB    6e38    1780dU'�a7�{Ǩ�Dh{d�����w�t\�J*��)���/*
���W�����m	��ĦQA\�Lr�q؅�fe�-I�詇��	���5�D̡R�D�88��~°v��]��\$:������FC�� ��>���G��;��в%z��ϧ�%�.�`�7�&�V�ZI�� �܈�f��U&�a	�A�XP�'�;�1m_w}-R��=A�bU�U�]ͫ¯}ioik;���X�{dX���?�)��Q
R�/%��34��s�S%�����Js�G��Fc;��?O�W�*��MC_^F�	�
�r�p�[�	`f9"3���粍�#%`B 8��򐽝r	v�x�}�:�)�a�]⿧_�=��HlGt9�vN�@f�� ��� >}�݃3����5�
,�����t<���v���X��Y�w�{���mbDNf�@���ϪW d�`������Mo�VW*��҈�C��	��I�8��P/Xᷯ��v�@���ld��� �v���xg���O-�x�ڳ&� �U^J%� �O3��}��<��K�_)��sQ�n�ȧ�r���]���Pe�� �nv�0���k����D�I˟|�<���%r�>�@Y̨^��,��ܳc��I�G�V_��j|� $)X��u��*I��?����g�-�#
 �+mH���O�~�6s�F��~��a����X���.NK����S���gG�b��Y�`5��lWBC���e���Y��c�	3��u0�Uƻ�w�6�y��ٟ �͉h�!��ĕ�����T�JH�n��3���$��c���И5BƔHb�o�iGͰ�MB�xu_a���<�>?�!N�;R�2k$����$�����K�~�+4tЧ�8�ޫ���-H}`��jm�|Y3;a���#GwC
��2xQ�M��c�/9�T�bѦm���q�����68e&��;�J�/a���B�<�"�����m�~��������魏R��YV�@�)�fi�#�E�����Ƭ?8�E=
�od���ߋ�>���%��0� V��b�8|g���i���W��c��R�!��Ҡ�j�^%䄺��7��+��ٚ$��h9 �F|����GrX���(�=,䒱h����"���l�=u��	PZ��R������ן˴Y#n���"��FN�X̃;�	^0��XP�b)f^�c_���������U4F�T�2c��keS_�Ϙ��__%�/h�!pz���#ra�o3Y��u�[�Wn��p�Z����k��|rM_���{9��p���^���2�%rIǜ��`��WPN{P:�L���+B^���)���i�@|횼���Sn��ˉ좥WT*�R�%t�0����>K_ۿӴ���G�� ���Ep����K��R*�]�# 4�i+j�FQH�_.����GД�.��1�B�ÿ_�_
9�_k�� q����a�o�e����K'dXo�������0�S�^��� ]9� ��x���G�W�
C�UGeP��g�t���F��==xbR/&!O�U���>'���QW=�`�"c֏;^~LE|ocR3�b��-Vha^Ʊ�zϽ�oV�f���B�����J��H�̎T�l�[V�� ����O��y�_��+T���������JTn!���x�|�mS�v��H��}L���^�x#z ��!�X�13���]��:d��r.L�T^��/�B����Z}���s�T�M�?���`�υj�f<<����vTm.0�˟]�~/]7#��t��"?������F���� ���뮯���vL��%99H���M�<D�$z��g�;��df9�eK:�i���P�IY$9Zwq/�h@�5�?o�\W3x�g�'h�X<�L�PTK
�$��c0̜�)ܘ�*NN>u�E��2W�Ht+d{�H>i_��l�)s���_�/1���u�dX68����m��Z?�.L�̜h ��S����z�X�Ehf���4n�2�
�TI�V 7N�!�2���z�)�J֒��fK$UP)��&��|V�?�[��x6)�ǹ�$^�����<cvq({��zX�(���_�����>��`��2��P���1&�6�8TN2��DF! r��>=^���Ő��x>ۼ�r����x�l�r��[6�G����� I�.ų�%%� ��":��ή_���V�ʰ�9���2�g@?&`a��h}�2����hol8��H��p@�i��P����.f�?J�	=y%/]���,�%�V�����j��Q�0�Ŀ(��/��}�_�\ҕ`2���r��o_&��+Y�cvJ�>L)��+�/p�`�nzkXէyB��3��f#�'�rBɥH�Y���2�X�o�jN8A����%-�&����n�l=��ȌVR;�����bs��2��58����r֡4��:65B9f��^=ɉ�GU�m��^��{ x����W��@���*�h��w�#}��������+`�2IW�M@��ܦ��
�7�Bf���$���Y���Cw�#��>l��f>��2� ���l�@q��+;ZAR������"3���d���ؒ#т4#�t>$��C]�,��Ū'i��f:���\l�
�z�lڞ8l<��w'U82mu�P�y�N)�~u0]1W:ޔO�1zL��f9�&�u�� 1!q�{��s��8�R��^�R9�d�[��`��c�|c�� zֺ�M9�:�^��5�ש�Y%�,����	F��.��Ԝ�������E�����=Sd8z��k�4`|}�Ûgdt�?f�^�p�~����	��ٝ���Jr�׮�h��x���CҲ��C�֭������"�6$69[�Hu�4bű��"����jE�<X��>
9Q�����{��~~d���7|�'�5�h����-x�����U��!�ƨm�]�f������{
Ir6F�����M?��~t�	����e���mϔ�*����;c�_
b�g���+ڢ��J	��I����?uhݬ��V4i
���hA�3{������s��*�g߅�|G����D��;��5 }-�j����v�����Ph�x��Bh%2��GC�K͞��xc��A�PG����f��Ұ���S����
�yΚ���rxqjO��ym���v��tȨQ��ۏ�ɑ���GC��J�3��nn�&��I�vtaX�-�K�����ۍ3��Vb�����[?��D7�D"um^�cmd���؋�a���Ŷ~����:��
C*l�TYܴհ��:�S*���|vʛT��2��N(zz|0?�d2���E�r�_� 3|k��z�'F�MQ�E��[��!�!��X�f >�ÔG��OY"~Kw���MHRw=�o�����t9@�er�Ӑ�HB,Z៮���u,�n5qC�=�%^����chto�N�g�E�F	���0
���U"D�5���*�k?p�g6�d-9픦��1 ��<^���Ҡ��2,��e��+)w_��(��&V[��x�o��Z@�%��A���3�&\R�ۚ�	r)��OahX�Scz��P�j_�u �H���5J�FL���Hf�����a�~L60�9��\\[9��u����;��nUT7=�7Z/�ቼט�ش�K?�W$^y�0�2�
8�GM�6��V��A�O���Eؑ1}.�g86�Q����t�eL�?
c�m��}��j��6��m���נ��Ug�+��,��{���Cm��L�6��R�܁ӹ妸N�+I�)|�f����/]qj�[�{	5=��)�ބ�-:��>����W�~+��$B������W�,�q������~.J�X��q�@�mة�}h]�:�Y�lw�y�k�D:��%��M���2�u6nf�Oզ�V��W�Hȩ����m�L�O[[��T�$ҟ�À������=]s��iҼXg�H/Ѓ$C~F�]Zbp<=2�7�Ԛt_��9a�J�Qu��˚�@v�%sfǍ!)����Nn��VS����{�Y{��2v����miI��X؟���p�ڸ�ɫ�H��P�E�
)/3/G՗��?��,d����f&��������Nx���EԔ�>[�Β<N�+�h��<u\G�@3�P�zI���]�u��q�7�-��֊nŁ|K�k>w�"2�<�l�Y4F%93�L=�D�ON�bb�N���^�����w?�8�=~�ќ�#Ԟc�ߎ�]�ō#�0�/?��G9�y�/a�������K��b*���!�t&3sT�r(K��)��2݌�U�O��Dd�����IѮB��.�o���$x�$0���*�ɡĚ"���5�.�(���L����s�px�~ ���|K��<ؗeV�%�B�!�qxݝ^�E��Q[�Ep&&�+��@<�-S*~{�Ĵj� /��BZw��8�����|�ԫ0ĺ��Z����1��A���BY��8�� ��1j�c*Y9����~���t'9�����w��ڕ t�G��)DRڶ�,�7��}B M(3=�fUZ(İMǟts]�}�����A�y޽~�����a8f4�mf�s�Kc��e�)�yT�r��=Ӭ���� �������r�$��ݢ�rz��>���nksj���@��q�jS,��oxnn	�X��T�t��Cb���G@���g(fT^1��9�;�92��
�U�eW?�q�Kj�'IU���q������{3���9$�� ���K�	��*O��tؠ��p��l���JdNV��u9HR��:$�-��K$C��0�ӊ2Ж�ԝQ�b�����X4f�l>�W�9��?��^曺��Հ�2�S�ty�i��,^L�l&?:=rWY��n��!�dn���ͩ����`�V6�M�a��-���ރ��4�q�r�0z�$��F�����~�j��&^~+�A{�w�=i&��g���Ⰰ8n�l��l����m<9i�C��ވ81o�~��	-���p�R�4�ý?]��^/����QX�]ģ����_�V����c����A��8�GS�I?�W�oQ��;�%��R��`�����c��b�7��
a�ǑYA�_LY1��g����P��Z��~�F�N;��Pm�uJ�����M��V;l��������f�t'�#�oj4���6n��A�Ku_�_n�ȃ��ƣ�ok9��oC(���۪;�c�k|#W&�^��hQ����Q���0���I�:c�/c�O.j����L}��S���6�P*��f�"�[��#3���N��i���Y�ڂ��;���v&��B��9#���«��Q���8�s�uRj�B�0Jǚ9Y �{�qs���`����G��Á� ��}?%�jz�3:0����9�g���l�<����}�&����
���cM�O���{���*�a�����s��qU4�G�AX�HR�ʶ�*�L�&�@Tϓ�x,�Q���ҭy)��+!��XcQC����E����@�?�׍�z~i�g�;�O����_����u��;*���(��d')vf\��`3�H�Jx�!u�Ϧ����3Ǥ����;��-�a�5,Ï)�I�D�ȩ�	|a�^��w��8�u�(��'(�2�N��s-r�V�|��0�|Ȅ���/�p#Q��/�\A�z⒁IT��4O	�"nA�W�r�.K!=�At�]�Ч<�.�E�'�Ĵ�.�׶�o/[R�op�P��V�+��VȺ��f�9��oOi�i�:Y%�Sb�����K�a��RE��A��M���^d�qAL#���9��ر�!�P���q��l�-��,4E9ɸN9JhDd��JQA�X�iK�U�A]WB���,��|)���:� �ay��*���cOI'�y\fNA�^�|���7N'[������b�d붹�RN�F��x�ۄx�R��C��1R��Eu=OB�	6̛�6��t̸ 