XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4��<�콅*����	Cc���m��z?���En�G�}�)�ɾϠ��[_K�n�/��Q��,���~֡��_�����X||
�����[֧¦q��\t~�5؋?�Y����ð��P�O_A��NN��X�+�`�&)�`�ȂGU�_�:��+`n��|g���W\�~Cb/5����t9-\��.u=��{�:��֥�η_�fT�ͷ�%M ��:vk� l���y�AACf4��7�b�-��xc�Ԃ�0����y���}O���?cW��`�b�f�c�MC�՝���t
�z�svo�[�A�Y�L�r���Ԍ�Yx����*�(mT�2�!wC�ltx�-�b���+�m��� �!��PM|K�s5�5�G{��ˀ�f�����$����Qul�|�����e��u�@FW�MRs���j`�u9~-kת˃<X����Qào��-DSH6��MRb��^�1�Yv��}�f.��5�K���%j�����7X�p ���&�(;͒�7�e�l��jS����Ro�����,S�[f�x�
�F� k��9�W�3��T޹f�$�&�+��[j�KYi�oJ��E�%�PB��"bI3[Q�Lw.ґXH�:����"��ᵻ'�����QN9����z�.�v7&0M�=�yu��)r?v,3ʮ����9��D�U��>lcc��a=�����j09S�E���z��_���e��z�y�S�3~Q����=o�ZVL�Ɔ��#�ɲ��!m�
� ���'�XlxVHYEB    4728    1360w���V��tT� ~N� c��s�����a������,ʚۧ���@�?3O��Ua��|�K�M:�S���k�J����:�r4��,��SISЊ��P�?��9QAvr	V4��/�+Gbw�<�l�ݚH(9	ؘ������j2��CkMkOZe�1����U�uƬR.c����PI�EI��Jk>��r=�*m�䗬�A��)p�c��hh�����u6h�/%!�[T'qw$�y9HG
m�A�wޢ��9�!�����WW-�5�Y 2!S�h�Q_Þ��T�=�����0��l���"��J��� ���Lj�&�<-��.4Y��O�Hl��ӑ����;�H�*t��x���f��`0�l�|N���~�!_����+s�1CQ���-b���9�þY/�W�<r)G!�!�{O�KnL�^k�%.�0^f�X9�)�3τ(J0y�O4x#�`�9+�%51�ma�MN2ږ
�tcLSa�, ��X��sҔ�|�kK \^}��]�dz �	,%�K���ݴ�N�^�x�(l�T�v����E�"}F+��d��0\P�;	�>�cc�L>Ow�_-��Q@ұ��d���=��QY��=S��@/Q�q�9n���!It��Go��c&~���qV:�DN��q~B��W��1&����`�C���LY�49AAC�\;g+� d�9�ʈP�,��V	��g��} ��lb_Y
Y������0m
�N߈�����ఽ�{F�����*�3i�R���1� B �'PO�Tng�2ke�L?��EE�*ɵmS�_���=ޢN".K��� �;�D���k`���"_��ӷ�x�RL[L~�C\q�����{7��.��b��tw_Ӳ8�1�-3�u���A�JC���8h.�?M�^1H[B�ed�d5N=7
�˴����E��=ez�a�w�*|���9�l0���n���o��^w�nx���b�����Zh���G8[z? �𹯄0���p���,�ɻ��=��y#d�am�$�AX���F��Xe�,��օ�P�"2�c�I�%��bJB8��B�j���͸���y�/��fw�����
�2Sx;�e��?����X����&���B����������`����d~M�/~H@��aq�st57��!�m&�A��W2a�J ���4�@�Ԋ
�)S槀��ǕT&�lI��G:�(��d�Q�
�&�NQ�˥̐A)���J��~}|���2�1tT���0u&��G���D�� �K�3.�����BR�a��vo�,}�d����՗Xk��6�2���f�	��D�`�(�'�/?v�H���%Qg������H#?�&����yl��Y���8��U2�J_A��7��W�'l��H[��u�]��te.;)�W�,�������ȹh9&�x�oX�	E��!��&�i�~Ӿ���d<�3�2��T���&;�~����Zi�����,J{CKlJ��C5e�!#"͇�_x���s����58����S3"j^%��Tz��!Gjs�;H޵��BfL��pi@XT�Ԝ�l��Z���w���������R6B�@	��oH���
�}3�6�l0���hDrx�gi$�CSJ�v���>k�#�u�%<��8�����b�RY�|�ڳf�� �`jK�u_���V(��ݒ�_���_&-2dg���OBeL)o����-�)��B����c�����ޛЈũ4_j��͉����ĩ����bov'��6A��/���(��-��
T�)Ɠ*e��+e���x��M�������*k��	���ROH�;���S����/�� J�}i�@3Q�o�.��6�A>cR
�r9 9�~%:�E���oN�)���Á�C�?�p/(�agׄ뷁�t�����^�Q��3f�[�qo���&�O�4Q�n�Q�d�/L�*�q�0ϯ��:��B�*���x44�T��+����" z¤C2rm~�ƋD1P���Y���fg�Zbm�B)��zg�N�6��c�K�c�]���� ri>pV��&��A�k٪�1
���ږW/QM��6v.�'ÀP��7��j�HXM���b���3=VA�Α�V������i3���a��A:(��oƭ�����_�_:�'����\���O����\6	�9��ġI�ɚ��YlO[��ԆG����̈\B/��ZQ�{����({��7�Y���T��׏?����9�̲l��ϣH�q݇/����f�|L�A-v�(Z�L��c���3)N��9�}�o6LKH5�O|�i����EF�%a� �AzIó��o�$�\T\'w��~��jw +�;����=R>�1JKʆ��VKz�ēg��^��"Bsw�}U���!F]���)\��|����E
sh������ȉ3D�������ͽ�����T-����K�&�]�l)Cag�#���ƭ�@�RF��8��%��&��g~��変�W�4A�l�$���>Ⱥ�3��B�n0A�Y�5fP�i�÷����[���MS��j����HS��S@4�b�ŕOes�݁@},{��U�b&�f����]b��$^�vWR�G8jؖ�=�|�D���q6����E�8���{#k�����փS�}Z��f���9"�\%)���q��,( ���x�w/��n����4�(�s�	HT���uWǎPf�C�����~�r6��d���	֟�w��U|	\V#���ǟ*{�����$��
^�W����i墛(PI����7�(@�֜0��Y���N��9bQ�!�@�`��5yi�,��)0�����s1bv�O�zj��m߄��/�r���
jck�r�*5R�v`�ƛ�}ޑI$Oa�SX�5N�R)���ъAE}���!)�%�l�"w� q.�I���.g��:��G��� >�P�6h�zz5'���N���]ׇ\����%AXrYB����5�����2ʠ���z�����GI/ߛ�:�������U�<6h3.��r�s�L�V��j�n
[�6��!zkbkz_��S`��q}G����Yg�3��j�_�a��X��Tq؜	vLh,!����_�$�FW�zU0�(Ό�E�b�41;�����9�S���
�������m��Ʉ�=��W6��"���b	7\ �I-;�Ы��
�@ʴJ�${M!T���r�tQ�D�=���R�'���MS�e�g0���z����+kZwVl#�<uvA�N*bM�`g�g뱽;���]��\$4�:O�r�ՉO�q���7ew��rww��h��0ChE�z�]9�h�Z=���ѢVB�={�Y��^��P��~�M<o�잆p�	 ~�Jk��Q�+�U�ڮw�2�Χ�l�k�D���/�֮.!�k|�x�7Q��b��]���2\
���T�y^�+xT�J�=���?l 1�9����ڲp�ft��D����f��`UTL���_b�0fߨ�͔y�7��/�g�ƾ(�ޒE�廴��<qN���`��\��nn���[�	�K�_J؞��Չ	�\`�NM'��:�Uwܺ��2U���M� �5�F��X"��X<�?�U��Q*����V��in&��K��j`�z
r%f����g��^��b�r�oS�Xy�Ռ<�͸'�ۚ�t��,��2b�7��-�R%{�#�W��H��T�O��2��J��z�Yo�#��H%R�ۉ]���k�vP\�,��!�Ȣ)��ϡ�GU	�A�k������-]2Y�o�0�*z��\ω"%��� �:�](��]r[{�tn5�r�od:Koi���rN�k5�2V�8f�	tj���{��*`w-��g�v��Ս��=�z�ߕ��Ej�N�����Y�֋�j��!��Y�55I~�|G�mLSI]��c)�W�I�L�>Ps�C�8mt��A���	lk�<@���ݞ)ש�4�H@7č���ә!�_ڳ�~]g���e�@S� ��E��V��c�w�N��#G/~�NO	����̣�jڍ��V�Ϣ\��k�/�+���~RlŽ�c��'���	':s�)��Z�"��)��ׇB�����hZtn�6<�+k}!�r���Ҵ6����z8�	� Q�ƌ���H�l:�N�ee��;߻I<
�$��V���+r�.sz~�@IC[l,M�9\�f,l�9�*�����{��|��S�T0����}��u�p��͋qⶺ �A�� ����<{�Z���mq�W����]2m%2�{.�=`��'���F��6�{��贪͒��bM�mq%�< ]ѱT�˞�[�M]>''�<d�Ҁ������䣙�n�L�L:Xm�+��ؑ}Xͤ�������G�˛�/���T1��j,9;�/��O�*�
-Տ� �;�h�`�&`���MA��k��CZ@����@��e?����.��k$��!e�����-^��D��T�NuҶ#��U�L��r>A�&X����{�k4�}T!��G�/�ߟUL���3��t�H.I֦��o=�^�o�ѡ�Q�d3�ˮS���8�H.m�~�ǃ�\�i���rKA�Y��UE�)G^`N���Dc�<Jq�A�I"�tăQ�_kE;l�úkO��K7>g-���@���&�_~�kA��Dk��M
��GW�J���<M���VK�>�<K�jվ�ꌺ�QU���[�pE(�i�?�1������'$be�����Vݒ�����U��ua�������~��t!����%@n#�ٮ�/�dU�Z��Y`���wh� FLWG��@k�Y��4N�KEv���8kQ�b�v��F/󏧤�W�,$��>�T'Y͙V�a��9�K��e�	#��	��s��w��X�8�g�^��iaG$%������8����5}�~�>i�!�؛'�A�ʶ�OC��