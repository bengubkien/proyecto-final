XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O�v��`��m<���{���!�}��>�8��P�&�`y��~"���N�I?yW�I�Q�{Ӎ�PH�&T�'�T��D��Wm���h1��ezK������&;�ѷ$S���W�La���=��2@z+��Y����|u� /-ڢɵ��q!���W���ס��](ɀ\�(Ǒ�Ў�q3�V(�R��ְM�6��9߱�V�IL��>x�8��)*���ip`= ��]�6^A�ٵ|޿2Gb|E���>9hF���M(��#���to)����f%Ʊj�'cQB�]�B���ݡ������	�� �+�9���]މ��{Dl�*tb�cme�Ƹ��&���ȉ�=�t���u������3 yhU�p�Qy�Vnv������o8*��� �fFo��Fj��$��Y��i$���W0�M6�USh�em�)�C����x��P��X�f�� �,2�����MrQáum}`��Qa(����ⱄ}�_�]s_x��+W�b��\3i�`�m�y�b��8:ڳM�"��X�ߵ��2g8���-0C�F�&VS�7�]@����f��`��|�|�����XtL���+T魑��i��Ѣ/�A�J5����8������J�\����oÆ��,��a9�wy�ݘT�NDJ&V&y����߼,��9����v(i�}����z�ɵ�����=�:������c�VkRi�z!_�S~�*5K�;i��|�r5���Rk����@ջ/�XlxVHYEB    1464     7c0�h*��#!?6�%_qe�����r/���������s�����b���5 Z�����A�1��_cT��3T*�3�����p;���@J�A�����閨F�Q�������<�L��M u�` ��.�2[=~׽�s� {�����ޞ&�E��2��ѶX�
8���(ˆ��i8~Y���)�}b�W���%�Z�7�,��;�W�����j��cG���Ә��R��ѯ0Zxʀia���*ֻH}�RJ�nE��n��N����2?A:�����%:V� �L"��U�	��?d�D&O�����]"xs&��O���KD�$%J6� �����(z"�������c�}������.�ל?�ukXO��8I��$�� >&$=��Y�ҖC�Z>�+�1�A�wb�i�ۄ����į����2�Jʞ���5���d&����|��:b��k̢���޼:r���ԝ�9�Nx�A��lq\�O�E����u���$�e�K�6Xs}4҃�?�O���GBg\j�9Ǆq7n.0�,E�F�A�ɩPw܃�d�V�=�o�
jYt��n�ݝ�`U�Z�i�)�h� �#y?i�XZ�f3C���p_T���	^Ҥ1��������^O��$���)�N=O���R��R;���O��tI��$���>�#�f�*��B�X���e)��׀�J����1��¯b�rE-��`K�w#?�������0��}/3r��'�f�r~:��r��V!��z�+��Kw��+���Z0��2�L*mp��q7�	�"ln��c�v����$	��vת^�� d�Ӧ-R�Vw�E�
&ȇ���Ԝ���Zc�3��jQLh���j'C鋃<uĬ](�=��
�Ml�Q�<p6�>��V㳑�3�C�j��ub���}Şz@�U��5�B��vEc�4�������N�j%��d�?@I���fJ�>�b�l����#���V��r�p=�7M����y&U����h���Uv-
�a,a�s>(3]��Y�VH|�ɟ���v�ҳDk�P��]%/��ikO��>�o�hxd�E+4�ۑ�p}��t۟V�#7b~c$�A��V<�N����t���ˉrL��p.�㬼����9�~ ��U������|�� �Z��P���Z%aΛ�/�vP���y��hr�>Q����'�,��������&��	��D*�l��yjX�'l.�HI��A�ᤀ�n���@�l1�>��I�,�h�7�.�)5���,����ҡƚ��I�\��7�3$F��E�N��w���Xm�P8a�@�	�F�o��Wv�~�X�;J�S�C��uP���"$`�@��+����Qa��Ёi����_d��g�Z�P��[0�x��ir�+�H-����z�?�eXW�Y&�s=��(y��j2���0v������N@���B�P٥l]ՉE.��A�H���j���Lλ���ȕ���~�[�r�^��5s��çd|��]����+��b�����T4�r���IQ,9|6���&�|۟�������A�\՗	)e?�m���chK��n�@x���F���?��_�r|^��s�إ�AB�a�"y���htI�O@���cv���0���<���a�	) ��|����,{RPp����� �M�N�� =��֐ye�ќ{|\(���֑m�=λP�B�m=�T9�{W�W.Շ�b�R��3�(:�~��Z��S��~��&�Qo�is-B�b�xd0_�����a
;�K�m��*��jԨS���\d'-y]��r�[�T3>��\C��ڝ��ͥ7�&�,�a��y/�-oC�c��4����
A�[�g�����O�PKD�a��nt���1E�����`K���1	�^�M�9d�(�)�@T��0�9�o�2F҉��n�*�^n�~�/�x�7�tr���JA�W��O����ڵ`��m�&�8��