XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��LQ�(lTR��Q�0�6`�u�o<�|o���ۂ�G��9�8$"/�a�ě�(<�g�f�����a�A0������ox�Y�>�Z	Bۇ�u��p��à����B��F�`���V�w�w�ԣ^M����Ŏ�YF5@K���P.�r���:!97�V���Ǫ]9��w��x�MGsy�T��D/��֦��o^(GH��#�3o`>>�\*VYN��b���սx3��Z�-UK�aJ`h=U�����_�O�jIzQ�eD���)��Y�j�<�Y����#��$�����kO]E;�?g��?�W����O�7�GT�u�d����>�^uV9�t��&��J8��b����a����@�)�!fPXoQ�lj�|y�Aw��<�j�	�g���z2�[��+F�=QVbX�v#�Ȯ�Ugp���{�dxx�-A/��@�M��+h�vhs������#�d¸�◇<-�S�?s�&A��8�����Φ����ݣF�{��G���X��m��V��r�R��8{��
�q�Ҿ	�'��}�Nׯ�Czc�qц�R )B�y�c�\VZ��ӂ�D���_,���P����$ɬ�,�zj����\��X7���R� �=$DI�$�* ����4,�P/�$�ALJ+�*�4Շs�t����U��8���o�2n��
~�*��U[c˧�z� �b�ZN+���,���P��չl�r}m������g	^^K~��'g;�1*<)8�2k����XlxVHYEB    153d     750Ι���SfA6^�s�Ҽ�T��A`!�j8���|~�'��k���¿K�5C���m/�Fp�e[����gz�D͍�-ϪD�,��P:�f��i��*9!\�s�Z��xogW)Џ*!Svu^.�Z7�d)u�-%7��.x&aI���e��~�,$[ �v����\Vu">�&4�K�o�O�I����Z!!?�]m���"�ބD2^%e!��tcB=3��|���銀$)�!I���.7��)��S�2���9����,�$�1�,��y��^�:�'���S��9xr.�ܽ����OҽkF�.d�v�^a1m��ۂ$�����RU[��W��jvG5-K�іc�5^����"Ϟi�r��L�B�{��;��%�`��J�tӡ8�	�`��yFN�߹�Qk�O�t������p��1,_��ȣ�o�'���(�m�������W�_{�:�{�K�����b%�\�� \�#''$O��_��7�e�Į}ܢF��C��F}�#��Z�!������"���oQ�O�dt	9t�!"���*�zjSY�%,��O�T�@e��d�Cr����WO��ߣS)�˙Gѭ[Tn�7Y�7��/��5��"�YV�l��m�����)�I�Vy�����mSjػ�H���6*$��������b�5�ݡ�p�5��)3>zG?>� j�>����x���v�e1O���<��;JUT�U��~�R.����^�.�_lHdC��]d֤�huܨX;*���Ӧ�f}di�٫��*��k~���g��Q����F�@�ޙ{тw�g�}a3�u���$hcg��I�l��&`b4�����҇��'k����<�dI��a&�n:���޼�߶6��N5Y�ä���`_���d>��պR�U��i�b�5�c��R��a�
Pq���7�f�Xoo��r�k�Uh�g����ޕ�R�T=D�zǌ.�ީ���8�W��/�B�$A$⍣��@[�e��)QŹ�R�rb��t�0^Ԣff-[��.��a�,`��Y&��2fJ�E'����X��(�u������۷^� PR*���*[^�Md�)��P�u
�齌��9����_�w{q�\�V��C��d	X�����a���GhSc�&�1Z"[$���t���ԌJ�-;����,�ާ�����y��cQ��*2���"T�C5����n/˂�^��^a�;�[�W�����q�b�E:�M�{�A��/�����~����%���k^~GśTň��d�'�Z����Д�)."����;�8�$�y�ԁ�V>���K�2��I�J�#��4!F�aʑpH`��a٧�����S�^G�_���������1��}�%�Z1p���W����A���PRR��k~'��^��θ~V���_�1�o)�KDJ�vm��#��B;�d=
�zJD�J���v@Hi�9yH�������@a�:�GmGo$G����t����>�G�� w���Er�B2��@��;>"�!|f�7�(v�a�C0Z�KP�*ze�*�B��^����ivYˁ��>U��eJy�x�V�Ɗ7 p>O/���'�:�7�cMܵ����8I,��:X	!#�_���C�V�uߵ;
�fϢ���lZh-iI2r�c�����~%W�"	%q�Q,0S	ϔ�2�ϕM6@��d4;�j8�S�l���kfK�)�'�� H�����|G��S)�@���r�#&i/~�r$�%ɋAx/o�N�������mY�n����M���J�}�0�W�����Y\�ґy@�l�Iσ@P�:.�3a�_�#,�Nd_s	J�|!d,�T�?�{X I+�H.�Dd��Y�