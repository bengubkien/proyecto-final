XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Kn�l��8�U&��ҽ����4�D�CqzB�:���>O|�=k��R��<n��DY���
�ʹ ��G�co6\St�T�i��q�<V�:	�Ԙ�ݥ
U����Ư���4,`��+��*�D�Ȧf@	5�\�*V~
���{�q�s!fv�2wa�$FV���I��l[PS�$�I.�v5���6���n����<�W����*w��i�g�[e#�9��v�������(����03Gx�ǋ����+�-��)�g���;�(n�}�ڟ�>M�]��������21�q��������<��j��L�&����޶��<q:3�j���O��k9=EN:���mx�``}��{���j9e�M������G��!h�cO$a� �g�,g0���r�6Ty���q4%��\��E"�kR$|�n�aYW���`�����L�����Q&�Z�#�t���JZ��i�'@�د��ޓB.4Iw�=1���+�d�oj��i��4�k(�'JN�Ћt�)��@~6j�L�-:�Ro���ԀF���Nt	rm$(������2���Ø�P���T(8�T���ZH�W	��D�5߃�%=��$8y l�&���4�j�Q���}�����(T��l���F���ES��GS�cP$������7#�V���	=*G���j
1�����z$�?m�T����*H���p�4�yt�9���wKV!YW�f��H9��J}��xU�h�r�
F�K:���$��r���XlxVHYEB    1b6d     9a0=��m�mV����;�Ƒ�@"���b��+(���%�K�����:R��>�����"Y�W��7ė��H~A��M��,�Kz�<��@� l�Z:���_ȯ�������;�Hצ�}�����\�TọQ5��	�O��A��3b֦2��8����H�V��ή>X��)z�2e��
+7�R���Ν_C�#�D��!�Pe�T����I9�7ճ'�5\�i��I����
���U�$\zk�-5y�����x��Q284@(f�A��5S�qذ'tJ}�$��d�zG	��EYk7�_�����\�C]��x�g�{|��YmcKL�w|�ޛ�an�z��L���I�Oj4C>&�*ø����π����n�z���g��0K`)wx�
��^2�"�Q˿�i�4��H��lm]Q��6�`����7B��}����Ɉ"7���w�QQw�7 ��!��1�G�91���l�G�B��ۀ�ʩ$��EbX�ؑs�Ի����� W.���<[�k��-bD��@Q^�� <P��;�_�	�Z�	��N����?����R���բp]��Q�y���5��
Ǿ�;��X�֖�(����[ɧc�HX�.����������4Շ��׬��-F��_/"'�����,4C8)� )��6�(�|�/�9�W	 �?���Rp�`�^��J8eP{|+��сr=�4�=L�7��]�C��&Qsf��,Lre�'�f+rY�����R�� ��ҁ��v����0����J���ؐ��������T/��C����Do����	�hͦ����/��h��!���gS���@�[��I��.n����y ��L�py����b�{N����\K:G�Z'��]�1��u`['^J%�v��|$������*�3_zX��t�eN�c�?<���^�3�[cH���9N�1*�O�f�<?>=r��7���
�qp���j�oGu��6bjg��d䏦�o�s�:[���k�8t����N�*k�!GT�_1�6�dQ��-z��6#��$a�8�<�4�ܩ�O�{����_&��)5Z�y=;#Y�2x��r"�d8"x��ƈKh6��<$�?��z�j�Of%�&����J�ϓ(C2m^I���P�AtG����Qr'-�f���E<���wa�S��� u���7r�r�G�!(����YZ�B���ى����m9Y3X�X�o�����n׉�<����\)I���Ȏ���{�t3ھut�� ���_��i�8�vj�C��/|��s���=�f��p�%Sϻ�l�� ��A��#��R��,�W �a'J6<�48�Dh�$_ı.x��݇�ǚ��VE���N�z�����q���ǛϤ�3��H��|"x\;х�
�t��辸	��-��~��������� �����k1p�A��C�	Չ%��X��:&m*:�`���J�p�}�%�o{>�vj�j�[��׀L�h���.�$'�������uo�_]�CI����(�<�R�ľ�N����s��Wj��_�;����K_��=���D��D!���<|�Y�n�I�d^!��B<a��G/�x����
�ߋ���(
�I~�`��U�M&"f�pu��qsi_"��+�Ję��9]���|@c�s�!�N8��4ҘӘ�B��jln�5��V�P�)�"�1�{����	巰��/�;dX@�A�	��>�K����2D��vO�t�X���zD����q����:����>sJ�&��}-�e�DJ�(�:��,�JW�|L9jZT�V$V���Q�)A��s��~8���Ԝ�kŰ��ew�f%���}�u���i^��]s�_��L���n�:�uB �|�s8y�^�{���#jl�ETs��,��n���r"-������{h��3]W<<��U�H��ʩ�{<`��سc�l��P�T��y���GrjT\p��U"�\�
�"���Y;��W��
�K��?��Aqq�p��Q�'��qQ��+�����'��w���"�#��3\uh|�܈���F��ݒ֎��{K�Y�r~B(ܠt'e�vt�n�Y���n}�v�(l�X��P�p�l�K�Jrݙ���;6���(�������M;�' �a�n�V�GC��C���6X	����-�@r�c	�e����jh���\����Ҫ��`��DI|�Z�;{'���
Q����fd�J��Ͼ7��/7k�E.��ī�\�v��Z�:�Uƶ��������G�iX�t���Ư��J�o=ߖ%8�C���BR:J�PD[�	F��+���䓞���ɵ	�28���&JDv���Ktu�^	��@�Y�S�X%<"{J�ZR����I���@���W���봯�?��y] E6�w�֝4%o9]|@�挽=����G����:0V��