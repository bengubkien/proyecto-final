XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o$F8�[K�ǀsy����.���<HЭ���O�'�#=UC:HNeƃ�$��6�d�P�xѮ���e/�S��͑����cr�X���r�q��c̿�݉�p�ݨJ�� ��Ki�RS��������c��u:�t�?��"���:�x�`���*�d܄�f`�V�ᵇ��=��t��j�yΈ�a�
f��%a�Ө�m�g�gx����{=C��'�S�p�w��K�ko�A�A^�#�+�VG�m�8��@�E͝�3�H3@՘k��1?��8�:�5z�F��>�P�cT{�M����w�¾2�dIc@����J�����j[��R��QL�?a!P-V�zQ��ǖ�U��hp6 �;�6�Hii�[Ů(�8N��p�	�N� ��\,=?���+<��?�Cì���[Y�,P�=��_�����7��(~�sWZ8I��o�C�Z��2����6ڷ�v�}!ͬ��o�T"� �O��Cӷ�1UsFE�g�����IcdZ��3�����ɡ�ϑ0:b�0-�������h�~`b�9%�MZv4�%?vlcπ�F`�"y�*K1�M���d����6'�#n���ӳ�:�^V��f{5Mt�c:���
���n�a�\��w�3l-��y��/KP8c��o�~�=�B�����|�k�B�H���(�p8��h�����(?�����HT�� v�a��/�iWX���4[�� �����2�w�^K|��j���ۢ�xƨ�V���C�DDg\ x|�^�� �X�멞��pXlxVHYEB    30f0     ba0��q=�X��cZ�χyIkU�K�n�E�(��.���p�<>�!�q�w}��� -�C�(����.��?��w�9y^�8��;c΃��i4�4d0��2Y��h��(yS֍��&�v5w(~��6��c`�7֪&��<�݌F�̯�¦y��{��&<\U[QoWU��� ��(��l������Aۮ_>q���b��?)1�.�aP�=R���S�d���%B�G,��|s_�p��o0��yK�ȥ�l�C����S�m:���������n*H�T�t�i��$=�(:/Ic!�wh�+?u}~����{�hm�g@�ћ!?k���݅ٓ��F��"��"\�/�S���3��xZ-q��UT��c����" ,g $���@��@Pw^���Hw��Y���H�4�CԵ	��|��zbZ+��$���ܢi�և�z���<�z�־Q�[�r�"�\�x^�Mr��''4��k��F���K���9����$*���9��旕&d��[��Vpu�}�A�Je9\��uiu@=~,<���,�o��SS�JQ'��� ��ĝ�q}� y[Ojͷ=����u�nBs�#;�W8;	~W� ��Ӭ�˥y#yK�� ��a�f$6O��k[@��-�u��0Zr2|]�D'�����.퀭$�!s���dy��^�'�����1tg�D�EAVڢb��Y7s�N6jw�����#��OsY,l���-??�z��{�X�P�����8�Ӫ[��1w���t�h�$�VB������*�>�I]��4!�N�L=/VK���..��R���&�=L���tf �d�;V���i%��#�z�Q���f�*r/�]Aމس~�+!w^�o�	����뷮
|��� ��(�����;^�$�4��o�=_8�d�؂7�f�N�Y��!��UqEZ)$������F�Sx�Ǒ]I9jJ]�O-g����v�yT���@"����y���V�G�pݏ�awh-\o�4 ���0��$�	�c�S�薁��=gG)mRgQ+W���tT��?[�jt]��|G��Qތ	U���
B���m;�xk�Ì���v3�����$�ۍRm�&���X�)���3�L��р��Q˸�0 ��u�723�ҧ�zkQ��>�.MWq��A��G@A5ċk�Z'�G�	����!�F81�^J�4��6�,Z�X�W��P25�0����<�V��*��)u�%LK���泝XvBX�~���\�Y+	�P8�������0^���o�+���B���⎲g�ͪ��(<2��S��74/ѐ y@�G��/��Z8��[� ���p$���}LͰ�P���7�4��i0�z~�,�{����j�um���^J�z�8��p���c�z����+NX��H�/{��b����aS[Qi�ȅ���ҐFdJZ� t�͗pD�0��E�Z)��0���o"�E�D����%����7�7jʛg�%^�nPpH�7�KG�ty2�nGh5i�[
o5��oR��]l��CMT����W�h�r̡�e�#��a���~��]<,�,��u �f�d.���Þ[�-_�^��K%�����c}�Q��q�@�C��pμ?��lG������&/}����v�b6ԥ�_ti�m���u��H�x��YF��WN{���%�T�r��kQ��
��c�[��s"�f�?c_���
�Lu�?ٕ���-�6�p�B{O��U����k��u�ٸu��@���@x��>P�l�DA~_�.��h(�k�֣�[ 8�?��;�.@�cp��"�p$��*��[�޼�����e5�y��v�ǟ�%AYF���׻kwk��\o�,��٪�#�2(�~�E]WL�����U�A�D8_���i˒�,~�� �c��������/^��/.����1��o�VfS�Z@k-�c���[��-:�ĐA*�FhU4V�)I�wL��!�"1�\yǎVA,E������$���)�
P������=ړ&�͒���W��o$��V�cW9r�W�ܷ�8�����!�GF��|3Z������ �FL﷽�</�}m�����)|K{Q�
4��%�5�ظ���*�A�k��oH�D�h]�k���Iw��q�@����=�O	1��`}�@��V�c���)�  �`�#�2�V"��Ɏ���Xֱ�N(#'��Y�]�E�Ň$;Z2�vu���'�p��Z[�R�3��9�Sf�7ͤ
��=Py��b�}�=[B��(�;Ԋ�d�U�/DO>	���C";J�m�g3{uz��W�&��h&SjH<N�Y�ʵ��Ҩg����X�1��� ����BI��6U�|%�bV�><��\�
A��$Ƚ�D_?[@g������'��X�q`|Eɚ��&���=FR9b�8je�oL�h��ŏ��b��b�!dI�!��T㫥�sV��^�5z�bO����۞����M��g|�(XI3��W�gd���Np�py3�5�hl�B�4,p��P�#�/AZ3��kQ 4<"-��w����?�$��G�rx���C�sX8&���ǶU2��`��-�e��ߨN�TÁK4m}>(w���������ofvx�,!�l"�@���Mj�F?9z��!�=ҟŷ:k
�w�j�i��{���� ���˝@�.��FO�� ��F��:����f�y9��pYK�������f��+'��~T���c���Π���<x�o�?Zlކ�j#{$�4�n��ߐ�T�B}g�A������^����.���%g�{�˥9P�7���r�ů ,nn.�[-4����Ù�T�R�v�6��I#6��m�.��,�m�]i�3�]��VV ~��*O�eG��8��f-ͤ�?�����R[C[_�PD7�HX�7����bRn!82���