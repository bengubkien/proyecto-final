XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D������Bȫ�L�8����`H=����ǫ~��lY!�f�$6"~�����/��E?��Qg1�zG�i����81Z/"�,u45�1���5�\.o�lxj���Z�M�i9�HH��J�yf���؁!Y��be�*�4��I0�־x���r��ƲIk�D'�4�O+[���G���xM..P�I��S�i�����Id�NH!�o�%�>�ۮ�O�%�o� �W�d~�N�BҌ�j0���J� ��͏H�)�۹��M��,x��VIm[Z�������9�4��q!fO2��1����(�:v�UY6��¾�<j�v	Eɋ�I����ݑa{Ak7��Xĩb�`q���I�;�x�E#���!e���֦��:�x�KB���@v�㟨���D���?���ʬaA���T7m�a�;�tyQPU<��G��$��14!\�55y[T��Z�p��ŷ�� L��DY��0ٷ�B5�ԓ[�ɖ�~^�b��[ʦ94vw�^��q��I�ρ��!ߗu�+6m�����0��:�VZ��d�����qw��,�������Ԭ1Yeͬ$��p���O��O�w�Ӿ=����B� 6�?�pMB���m�V�og{��@��o뺌3����,ʚ�W��c/i��b����5�F>�C��Z!�&��Gٓ�.w�h�CQ��pxfW�oO=؛�G�{�����������i\�Fy�5d����׫��xu��Q]�Ǖ�g��i�m�>���h���?+XlxVHYEB    2fce     cb0�@T�Մ�z�`�	8u�ā��-��yz�� H�Mk���.l3�����P�)�����S���fԤ�f��h�~�,�M�+4��֞O퉮/��\x�rE������]�Ԧ���'� ��˼!���a~c��/����@��?��`���'�����:�.�8��n{���,ɢ�Gn�;R��ĵ�=߄��b\f��X��EuE���F%��\�`;�M�����WRg��Q�����]ڡ&]P�d^R\��W�������a�q�	�{�q'5�쟀�xѤ����n_�}.�_�N_T����J�{�]l��
�P�i6Vz�������G�t�	'kr������E?gq�7�5=:�/�[B:�� �,�Ӂ��"9����L��S��M %g�Ť�*�TP����?��򈈋Vp���Y���p�w� v���l���y�p'���mN݈�׀R>p^�;���}�tG�j/� ��	������S��À���j&s?j�qp�I�v!+�񫘄�Yu3]����y�.�pk2\	�7�f��C�Qu4��� �\~.r�De��G��]ѻ]�1�D�����{�d�d?o�Opӛ�"δH���Bo�9�/����,���HPܪ�p����x�]h�٩[��D���}��fm�炒���1m�(��A��X3�r������G嶖l`��&U��X�~�	����F/����h~��7��0�T_.� �-KZ!0_�Sc�9���5Jмg�:����J�PǑ�˜��'?O.�����ׂR�@d��kl�!��7.����?Q��7�P#�BG@�"�>l�1���^l)�U^���rF��cC� %��:���J1�T?)Ў��0߯$��=�gA��A��,���	Y6�dɋ�{(�n�Lr�U\���� D-IF�ܛCg��p(msY����"<�[�1P���?� #_F��^�/��4$���%m��!���m8GT�S���A8�'���2��h���T���V����o�"���ew�Lg!����g�]�E�
��3��_��*6K*1�6n*��U���\3���*s���i1^��	���sZ��9�xYц��p�i��m��ނ�L�\P��UO�g_��Íp���_hT�ĈA�Pl�99b1��jGL��n�ԯ�ց`����%ӌ-;��7��au��ɶ��֗n�[ {uv~� ���f� �*	��f���
�Q��<p0������B0�(�E���=��C+C��Fc�=0�&�k'x� +��U������&z#!evCG0���J��;��ǀ�N�~�w`��In��P�6&;+�Rb�TM�ѭ2�%E�{�U"�����A����"5L�ιԠ���GYkE��'��	��;9q�./N�@�*{k��2���������w�^�LA�|����ȃ��W��ѝ�j��;;� !�M�";���"����FKp��Sെ��oH ��H��=ǧ+W�5*gf�����Y���cRJcQ3p��C���F	m����[��D*v �+���e����KN)�z��*Y+{5q�[��]��~�5ڸ���iqNr��ꪲ�IE��t:&	���pܼ�gZ?Rԥ�E{?�d�.��#�K��<h�н��dcߡ=��5Su*RL�^��;�A4�Dۊa�q��s�o�39�����н�w�2�,��=�L'u JН!�'�}���&'$�t�&Gww����a��YhY.Z�i�,}�����J�)/��+FB�j��X.�*LеcK��KL4~����b�����v���-n�ZP�e�z�Kz�8��9T�dv���M����SH� -�xؿ��f���:��rv�ڹݍ)��T9-Eb���*RL��܀[.�O6��s+G���<�2��4�~�>B��m�+H�i���;ĿS[���-vwz��n����@��0�7ɋ������,Ǣ�b�j��W�	���ۡKh��DJ���`�Y��;�P%�D�47���Qe�̾X���^E��7S��"�2����уW#�(c�~
]IWQ��fY�lMA���#"a�ͬ9ƌV��U�Њ�|�fc�*c6��Xն�t�Y�������і��q�� ���@�`����M҉"���Y'v�gl�c����:��s���_���� ���[��o�y�;ܼ/��Y�4�YE��>���/E츬���e2|�zڀ&�NT-��{̉�J�ޛre��̻������Y����G(l�]�8�ݳ�}Ӟ� 	��>uw: `^?�����2�`��y��fb�ˆ�V�$�k��p�Z,�Q��),�_����t�v�=��慒�u��){��n�6���?1�\�gM�K\�&�eo_�Tx��n<��*+��Zq�V];��	}�`�� �.��/��x^��7!�p��o�_�IƧ��s"C�̈�`��g�Nԓ�/��{�?�}���!$w��/�bd��~L��a蕤l��}�pg��{?h���o�1�����h�������.�YN�U�**�q��?2/�+�v�L_Bu��='�����{4V�R[�%�Y�������GZ!_J9�/pBxb!�`�N@z3��Љ��ӻI���\d�l|��M�P��XV��t5�����t�m�bAbv֥��d����1q�Br�zl��'�,��FR�2%�U1��Tk���)z,�α����{�b��u�`pvyu�z܃<���T��R̗���視\B;?�mPg�{���۲��T�D�������z��H#�䰥���
P
�j�oռn�q��<f'���{?��N������KA��O�͡L���Շfj����E��?SS������.hd;pv'�}�{3��M�/��̸��=Wrk޿�R�+��/�	�y4!�z��,0����bZ@NՂ6��25];Vs��L�u �9U�'�o��fLQ>S^������S_x�.��я�@(�sw.Hf☾�Pt]o��1�M[2|�6&�nE ����*�@����X������8�aS�����`ɟ7�
� rn S`��?����ܯ��?L]B������fO�в��vN���Ծ:h��i�_[�e���:�j��I��-V Z)M84Q#�n��M<ű�+vv5q�DܲF��ѹ�U�_��Kd