XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s 2�|�!�)���F�=�x6@mg͓�+�
U�V$A�N�r��Y�j�jld�}�@4kY���)�\A��*�ݶ���O�q=s���)��9�b����-�T��e��jNR]�Ģ��	I�6��%"o19F5�'�'ĵ����F��
�-x�تg TxuT���/Ū�Ӄ\�F��z5� E�Q�G��Amt��[�{��Ƒ#�R�G��ܧ�/�I�9gA�$U�_���T�F8�_�,�"�������~�v��Qh�8�%٥���<���ˉI�/�������p�Z!56���/U�yI��:@ﭱ�c�5��C��T�9��x\�uU�!k (,��*��'�[TU�q�Nl��qޅz�B��	�A�.��S�{�ɀם�#��{Vr�K�Rn��,�z�b��赵M��Q��&T8��I`���I�U %��3�(�����L[��_b>MX��M�����b;cO���3�}b(�!04��S�#�*?���l{ő>�	�(c�O�z�BM;�����)���c�AI��Nݮ��I'�!�>�qLFc3�Mu?14�H`�+Ǐ$2�7��~a|���c�Ak;RȻI��!���ø�B�F�]���T�>=W���K��zux�,ty�L4u`(�gJWi�x'U٫��n�����
H����{�9Ht�9?#`�(b��!�
� <U�s[�"���W���(a�6��Q-ܗ��,��	J�����|�,S����/Q8xK3����s t{���r��XlxVHYEB    6511    16d0�r{,u�bn
E��vit�Id$���<%�<�*Ld���õ��R�n��=M���k���)S�/���l{9ZCc��ne�1��D^u �Q@r0���`A:��x(]�̀���D�)�� ��^��~�+�h&���;��`�"87��"�i0+<`���;��+���� ��W��j�0(JW]�MLf����.j�VC+�T��x>H7�<�@AaћF�C�A�o�m�(�9���\�5�a����fM%RYV�G��^�d�\CfZ{�&1�d_�݃W-�V�����1$��H5��;��T!dK�;ڑv,"����لK��fz�L�&`��}~�GD�YG�[�4|��a1P�U�!��kK���Xˠ�#�=d@R5��K�4��[���R�+�*o��;x�R��^�X�8��j5��L>XoL Թ��]m}#[�=>��>��(s>o���]�T�5J��B�R���W?�<;�)��	 ,q1�E��
��N N&��k�cc��>֤��8���V1A>W��]G{���-�f$9�Ef��(8���+W6��'[���[�D|�@�{�c��<I�-����P�0)Y�k�>6��ۅY���t8�Ԙ]?���^m�8�jh܊�p�N���r���iM#[ƴ��{:�ᔢ�o�Yqy�5� ��
�ׯu�U�~P�^/+��ş^�#�˂��m���+��ʭJ�� �Y�(������ҙn-+���D{��(���a��w���_�I��؍|!��	�13����9���L~; �����g'�P�3���#o�i�Jqd!u�C��xֈ��>�u�����f��ˤ��fY�-&�Hv���#(CؕFd<�E��q�k3v����N��1����^SX��+ڴg`��H>��R���س�/����Ĭ��F��Y�8�U���S�o��!�-Z��\!�)h�����Y���=]v4g;dB#��ɛ�f B�IȆ.��	���k�5�"�0�ԯ�����T,�q��^���Eڹ�7~�j��Ο#T�Y��;%�8=��j�,?����ˬ_� �?�X?���)'��W2G�"��Ăoڿ�%6�E��\�9'�%�;.%�unVn�F�&���g�C
L� ӯ�l�]q��c-t[�Xc�]Z����[8�W���[�킌=�|v�t7Z�����m�	J�JP�N�*�=}ď,P�G~�����ϔ&N�[�o����ow��y�'�Յ	Sg���d(�AS�	�"%�.��"��Ϯ�pT*^m{��v>�E�դ�M	\���[�i0y��ǧ�h/������9 ۹���rW��:��f�Rt�����L.����4����!��;w�5]6<D���[�������U�x��KL���ӡE�e���Z���5��6膼P<�C�K˻���U��c�jZ�eu-mzyjdXD��fۓ�p��l��~^r{�ƿ�����(S!�Ew��`�!2���:C��(=�.jg`H�Q>7Hs�Y�����<4SmU��������}u�~8�f�d�0�mG�Þ�g4��.�{�%�U�ꖉr�^Gpm��/�dE����3��yPB�8;\�.cO<��3������K��D������n]�f}dy�{�Հ]���
�/E���E,�3~�R��LM@m&�9��<ƽ���P�q\�r�^��)v4�$�^�/�f�7K<�����zD�z/q���3D�Ν�3�Ձ��/��*�M��v%��9_�ƴ���b�a�\��鹼?���=�c6Hˇ��贾-�T	HVf&���9V�#�WG`E�&Y����l�����yh�rT`�S����̝����f��p�'��r��
��`|C��Am�P���h�T� �F�>�J`���h�N��dz��I�ӮgN�p_.Lc#'�ܣb!-��ϔ�?Y+�.���:���m��Q1M�N�]h�KɎN]�� B�����MλT��I�#��d�1\1N��A�M�/�_�*��B��rVm�$ml{��Uj5�Q>y)�Qz� l�U:��8ܳ\"���f�%M󅠍Id;���&�������6�����A��5�d���L�M�$Wd�R�i���6���:��ɸK��K�sL�X���w�Be��w���b$GAzq���^ύ�E�,4DL����
�
��a�s	k	���cs�u�gн����{�@���R!�.�RS��J��ÈW� ����,�vϗ����]D浚����M�H��ۤ&�ަo�V��=�ڔk7 D��Cd�Y�aC��� 7!����T�Q���.X�������0�Ef
&f������<�zc6枠L� ��4��L;�	��H�2���(�LÏ��#� '�
�*�!i61.)������g�I�X����P�IS�*2 �?b�wGz��}���2�
:�~���KZ?��(/�k�1�l�gvz5Y1J9n'� ��O7~�c/�g�͌7a�[<�\���;^�6�|�E�Q�,��k�р�h&;�M������h�p�Y��<e�s=c�9����V�3������g�`�&	҄�M���_+� @y�z���On��3]�z����F)X����J���F��� �g�Ve��G�mϖ�'�o�D��E�|S�u��m���:�&H�E���Oϴ=�F���*��Ѕ��ܷ�}ӢُcJ��	$6�^ac��'�I���Z0�/��Ŵ���<Hi>3fr!��}��]����)>�K�8H���JD܀��Ùy�w� *�T�@�511��1�I�$;e`C�o)%�C�FsJ�FQ�C�,�<Յ���!����7�~x��#�,g�<l/�2t��*%�<[΍�������X s�S�=:1C����a�a��}Bv�~'`8�ڮ���*��C�Kh�U�L�qq��b��QC7 2&�Ŕ�������hE�j9J��WeHI��22oA+W��s[<��D�D���z(Sq���f0��+N��х�8���k>(v�T=do^/�PǦ��"/̹��P��z6�	f�2!��z�\��F�j�"�pK�ܸus��A�Y���,@�?�V�;���y+0���*�RW�WM��<�����貊���LZ�1�w�������)5_gbK��=G/-RQG-/�����ӆMXە�'5�@ |
��M�Ս		���A �����R�F�o �\� :A��!�y�F�e�c��S���?���'�/�����{�&Q��M�/��3,�!E*�~>��Զ�
� �����-�͂� D���iLs��
�P�d�
�)�h����L����y`��D�*8c�.��3z^�D��U��:��@,���|Y���p���lu_̌�T�ۗ��Ҝ,-r�(1˳�}��՛䒖ˤ��K�}u������;p ���Wf.�h�-��ܧAj�,ÑZ���tǰ7Py��]08�k����L�z,0lh���w3$�n�b"��	�
��l	x�!F�.���q������K$��s�T8��ڀ��ˤD�%�
P��V���rtj�X^��KU^�����h08�6�a�A�jQ�7�a�+�� ��2	�2W�d;����K����f:�FI��Y�/�8��=�ԔݼK�;��P�����_2�_����U3]�7�s����r�ҳ[�V�'{v�}���h���/��T��?$6!�Nz�r&�M?#_�j2�){��.��=�[�	�03y�[͔�KB�I�ag��"�"M�G͝�͖�2t1,)$������PI�rC�\�w� ������Aa�f�*RyAa�äk}㾦|�����*93Q�m���ƼEqI���gm�#	*"���cA�����!��#�~]]�����Jc��L�5�$�h�]��G�4U�ܘ�9��x�S�{0�^�����3�3�+P��5�3����^��p����W�=��T˼�ݨq�cq>��j��N�l��/� (.iIA��	���vp.0�
Q�ɗ��Dq��L�yA�T֮)��Mz%��:�F^�a�//C����zS���٨�%Kl����,,-K�C��r2��ႂ~y�7�|�%	�'B���5W;x��rr4Nh��ø`a[fӢ"�����~�-f��͆opA�I;�!섳-���N@��iF@�j�)�G���T��Oo�	�#��ެ�>��o~-�0���wX�'���+ﲈKݾ�������0'Y�'��w��\?ԙC���N-*b�)�j��`<�d�����,����w]J�o~�8�z����{܀��x"��z�a�2�*��8��I����Y��m���R�i��
��G�X
�QP�En�~^�����݈?�G�u\�B��X�E�TY�-n�r�@��|��kb���:��2*wg ��<K4A�,�!�Z%�����P�bZ�tdũ/a�:�� �eO/��դ�jf,�7��j�IM�M1��b=h�p�|k������#�Ce��?|u�m�����U����Nn�o�v�h��vĚ8݅�+?��Bz͘-H�&�� ���TT#�WV|��w��E�x�ThGgvU/`L�6��/�:��8���������k��I��6T��XC��)�Y�VR�"� �:�yIk��}���`�8M�.�ô����-��$��4�c�i�EB\f	���쪝�#A��Wc�������jO��U{t�#�&����#�C�2|ZA���6�:	񺨐B�����d<��>��!p:����O�3�D���܋Ce��
[5=�?�#,%�v���N+���f��e
�+2��3�C@;��P4�����YS!yy�P;Le�y�&v������Ԗ�/����릞�g�4�C�ق'�n-"�{AĽAq=��m[��a�S�s#�g��M��Fv����f���
�O��W}?|��A�*0��Ez/�P��z��w���ۉ�z�d l�/���v�F~QN�r�$�^�{a�V��j�	V6�GR����P���<|	�bZ}f�Q�Z�\8�w����6}�fe;m�	!���]���=�-�x�?�����s1�]�r5��i�&�Qx�K���01Ltu9%��Ŕc��Ʌ��*PE�v��G	��Zf{"�e�e��؝A��|Ϊ��L���qk�VW����+�m$�������!�]�Z��jb����SH&i-شp�r�n���C�2	�h�<��LB��6��K�<VZ�SG��-=g�� 7ⴇ�sV΋��>�}iP�M�&џA)U�\ɵ8�pv෸�h���9?Ǯ���1.�M-�5�f��PS�!5��9E�Y+~5���Rϧ��|5i����E�NY�$�RR���	�U�1��Ѽ����-Go]��O���ig�|�og�21p�4�t��;���]�q�3�F͍��xd@zi@K�����'qg6�2(���m��_)�������:m��¥z/��I�-{0�~��&�\�	�E�U;�A��u�^�c�Q��i���v�K��M^�\&�p���DYj� 1�ސ{���[���)H�<1��X;�"SV��d�M!Ҟ*�V�~�vx7�	��y^'$iM��(���t3Ezv�8�� O�N_�(F~�;:r������3@c�Ag��A3(���_M-=y$XT�e \�Y=��������릁I<p����8ޔ�I��!?�ük"+�l�gp��+ ����K�ܚ�Ǎ!1%@%��y����=U