XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x`�5�5�Ճ����ۑ� �;�H(:/�>�Lj+�S;l� ��=U������iQ����rfuS�	=��.�-h�ϥS`B9v7�3>�Q6�5��8K���9��n�^���W�V�"��/�t�;hf���ڭD{�}Q���V�*N��<���R)�t�\z��'�2�H���ax׆�{qܪ�d@\�g!�Í�#_��i&=��9�	ᓃΊ��xF��T`zB͡]�I�<:�Ce��T�X��d*��t>`�!���	D��"����\�	}����8�&����CTle���	�ӣ����ECR�K	/�����I{�Ȭ�,C&�%��A]Ρ�Q��ˁ��� ��w������o�\Y�c�յ׀���Gd���ea����M%�	��1���H/��@;�S}A�T���g�^�(0F����I�H��H2�]k�9���"�^n뛟{��(~�������B��A˥Hk8�y���e)W�p��*EYF�����i�<'��&p����/b�U�?x�C�li�&^ś?I��ˉ�">y��N'�x��;�����6���x ��yPqg�i>ڬ:����.
�L=�|����5i,���1Nw��Tn��jk7HC��<@�9U*�Ӟ�T9�� �0�9�TWs�؟ZuoF*S^�4�[��B��*x���a�}x���&``������KDF�#�*{c#��bTd L<�H\��+�K���4(�̜a�<V����KӠ���:9/ѝ3XlxVHYEB    253a     d20r���Ō��]��˷<�p��-w��p:@>�~D���@�|��	��<n�;�jK�6 gh?�Y�Y���4��?X{2�N:�����?*���|}�O�����ث���C�-�	�
w��L�e�"b���Ό��|�B����Է�ΦlDp���/Q:bc`\� ���D
h_��2���<Gk��#y�'R-�3m�vdN��O�x P<g�7^A���1����0!Au���x �7���m�;3^�j��C�[FN�S�00K���n6i}7:;�����t<x�Lo������C��ۺ)<P�]3��B���\��'G-�&�6��ښeA�:/�5^��������^:���f�L�)vx/j:A��b12
lnr���ɠ�1���py�]�?��W��������x�y���-��D���!�gQCز3e��2���E_5�a���L�Ƒ�?��H8&2�(�Z��6���0��������|��>3�ҳ����l�!M��~��(�IN+	�(#s��Hh��y�Q�t���������c9�@+W�Υ�"���������&o���͚���b�|��9}�T�e��Պ��l2�j�/{���8�:@9]S��A�8Zr���y�1�|��w��hm!��Wȇ6�pv�xQ{Iۡ�*Тh��@L�̯K��1?&k�w@�Rs)�l}F���yo�F��E��u�".�DayrJ}��jq��;�İK㮳 z�F�-�mቯ����^3CQ�JK�d�sY��%��y��R�ɥ��hע�/,.m�#�Ӡ�"���Ϣ"h��� �P��]�Q�2]=�?/���C-�V��R�������������c0%t�����~���@�8͇C��]��B�4'���(��*��5(��G,���6V�.�_��?k�=��ER=ȋƔ�������]�ɯ��=G��O��-H�qG�/p��b�F��S:ܒ��PfԢI���Q景[�D`��D�2x�'d�R�L�𠳉�}J{�$B	���;����Ƃ�{��]�b����E���c�L�6nD��@����d��6�=H4Y 'O���f9)<Ш��`�\�Fw: V�1�M��@��b9b��{R�_���m�^�^��}�K5�2��iٌ<�	(�pMu��-`NRk�=��@�4�d�`�E��HΪ����&D�>���m5��wϨ�x��Y=$��O�<Y�A�Y���K`�(�٘����E�m*�`�'��8֩��O��P�Ԓ��4r'^
�=/j^��/�y�#�F�4�~1{J����_�i� ���7|+��k�2�%Ak�|�b��S\`R�]��/�z�"��Ϥ�7�N�k}���ډ��K��4|��GS��B3��; �n�r�s����u�������ʜZh(�ܑ�\� �bel�Y�80ρ@���*�Z�-�����qs]����73��
��3����l�g`!�w
a����9hf��5x�}9�]�����#���=S-��ul1�7u��f�KhM�"��D2V���wc��*n���fB�.�*tA����F�Ս���5Z-�T��HԲ7�2pxk����_��֏ �\���r���]]�Ռi�RQ4���ȁ�Kܤ��,ؐ�-��~6�I��q�4���=f�W��H{c�A\��}?�'M�;��Ő͊��$c�bxXf
^�g^�X��0Kwg�����eӧ#V�d{��'~���y���m��0�1��ӂ��))aq��ncZ�al罭F=l�2�9�m��:xd�yY:{+(0�|����@��j@a��/nOz��	�$���(5�����(TQ�-L��Wq(@�U;v�E\S���{g�:�����3��`��[�H����v��@���`A�sĸ���V��2&f%Ȯ�e�d�#q��1�U����=q �x���o�K�V3G�B��c�DI��赱d|8i����9z�[��_:�4���pxeiԦ](흱�@NQӾ��Q��Z�7x`�x���&�2_2�t<�������nd��떜=.�x��o~{:y��K�D�q�h<�(���q�+��@�U��NZ�9��g}�멁@�u�k3B�G�Ĵ@�tS�A�� {�%���-;�����\҇UKy'��!H�u�*��]b�k���V򶕇'�-�����S�W����G�,�?-��O �Yr!�����Z�	K�kB$4��m*v��*,$Q�)]��>���L��O)��U��o2S%i5P�#K��"����Vp|��?�6����&qV8��t��q��1��
�k��Al�4; ��ԩ0X1k�N�M�_�P\Ӌ��?7$�N�oYl:��NGS���-,urHγa?GI�[es�͓|��\�1u�g��`q�b6!�<��k��-���H��rv��)A$����f.n܁0�+�Z���e߳���A7)Ta�O+$Z)�Dϔ���Y�g��TU�?�������4��p+����L�I��|+�ׂ�1:�/�Z��N�s�t�X�P�"r˕]���g�8�Z���T*F�Jd���|A�K,�����ҟ�%���g=���i�1Y#$�}^_я@�g�/5-�!�σ~��TE�q�io���p�
+A�:� !zr�W}	��XF21����,�:��4�>�.������8�P�77"�g���(1|��4:�Bq�bE`â�f����E�V+	3搃�Ք�[v��D	��Jd6.�P~/����-Zn۔�8�E�����U�����k�Ƥ�B��b���g�CcQ'�>�M��W����`���g��'l��?�WT"@vY�ܱ"Zڗ�|w�&F�8�A���Gm�M %­T���F˶6�&��-�ڏ�a�Μ�BKY�;$��Ԭa�8Rxb0�Y}��;�
����lά:Z�ڊ8��_}L�U9��9�-���
z{��U�Y[?��f���WxJ��c���+�D��S��S�
�_�Ke�����������hF	��G�����A��s��,D��mN�k\G���K�s�'�?N��+D�sI�T:k_H<�� "�HK�#cF?����=�)�W�Ǽ�]T���}m��,Ǽ���x�ql��r��j
�s?�����iC�M�3Zu�Mg�ȍ�s��2&w�T��i"�ܱO�M5׫��d5�����#�|)�����P$����H�%�\���eV��t M�khw6Sy�&�.�
��^�`�l?�N�>��W��!r*�u�ͭ��d�`T��|�v��O��Z