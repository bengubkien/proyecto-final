XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�F��O���-Fu�O�Vf�#�ѱ�"�P��fꭃ
:��A�`	0,j��1��6CQi|}��j?��(h��8�)[�����Ǆl���J� ���r|���
BV	��<��@\�]�db+��#8K(xt��ʑ*rT�f��8����S_�fo�o�|b��^٩d���V
�r���	aܛ�T7�)�-��ƿ�JCi�=�4�u���.�����3q:Қ��ړέ��"�2j�Ҥ�Oz�mG8b8'W�	��<�\R��?lO���uY�|��sH/�O:Y��̥._�9I�pȣ�C(�r�`_ǀ!|>}�)#륃xkV��wL	2s[u��l�a�x�^{��	��n<R^�%5����CG���E�M�(��L���E�:t�%8�u�65�x�`8wGd���J��f�I�>��vrvGR�kBm��k`�zk=������ʼ���#*�);��[ �*,���	F��v��8csZb��f0 ��HA��p�8��I
%�0��18�o¸�a,&V��^����4GZz?b�
�u|�Y����3���^|�l���M�[�A�J� �
W�i8킕��KQ��SLt��~u�	%��zy�R�h���>��j=}ɘ��EY���P+��3G��xB��y_�������΅���z(C(�������"�!�c6f^�rտǁ~�-������A��`��S1qC<zafʦh�jc�4N�a7Ik���E�6�50䣅K�XlxVHYEB     c9a     610_�����}�QWſ����_Gg46���++S�Vʱ�U�)gbC�� �K�c;8TG��(�$�MR����"e��.�P���P�sf�=u��(�M'^�WJ���R�V)����`���͠�J�� а�r1J'�'���Z^��_T_���d ߧ���	� � .�����}��C{�f.������})T��6�C�k�ˆz�
�濏�'�^҆IY�)^a�K�\�k*� �n3�pjK��4��7���l�5�������i����ȳ�y�eK�d`��D'�b�l��DSe��m�+��x��W��cK�rx���]l������h�����~q1ƫo ���a���4�k�~x�?�:��X5r8Bygυc�J6%5�������nuh僶Oh��#���Uy@�� �Z�^K��1H�O7w ���`D���E�VF9(ۜ������d�1G\���&N��PhC��������K���&�{S	g6��n=ƴM�t��ːJ-�{S9���!����Hޜ�;Y�1؊��^:#��˰#K�㴢�gJ�2�A`�^�+8hsnc��l2*�$8�[���Z�{c��qi��&�9.�IX�y�N��rM��!��OD-��r��%�Ɵ�5$_�2'�Bv:����~r�du����q�ꓯ)2��yJ�g�4�5p����� p����s/�7���s3��b���Y$��CKXA�����n{㹠�Ͼ�ϊ�G�|]
�۝K�KC_qz�&��#��p��\>_eP�=,�s�tq�80zkL�'�b��8��<asQ���;l7�W�/��H�B��[��{��v�.���@r���B9�7ͷ����6�Ҥ����
��8_��ʆӿ�IV�����v�iS�K\�C����Cn,��!�ܦэҏ8InEe�|�>�,a!�kũd
�.}�;I��_�l=GM������E�2m�Q|��OE��&mh�tC�'T�O�C����x��������џ_��6���WO�L����nP��v��-�?q���ˮ7��Q���p��Y��R�,��{~���H������I3P�S�8ݧW�B���R'���(�����V%D�0S���)/��$J��+�	-����"��%��bs�<�Z��MHR~K�{�LfS��!gk��O�˷��	�r���h����0��!&�Z��ND�sWػ���MN'�c�`޳���d�>~7�G:����k�?�[�?�Q��gZ �T�r�� ?	ծ,6��H�O7���� A�NX5�v9�h�����jD�*Ϩ��nA�G�S�_D)�R�#�b�g�J��k��g6��d�g%�5T�c����DG,�h���1�E �7+%�eŀ#�������|�b�]�P���1z�Dȑk����ӛ�:�ZId�4k�@(
���bg�u���D��׏���}1��k�x	B�U JWE�xP�L�ݜ��N&�Mj�:u�KևƄ��Z��gs�A,������