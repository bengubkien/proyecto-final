XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��|�d��]_���MՊ �-s@��"�:�ǣ��ӕ}+�u�b��0������4��ߑѡ��O������mҚ�f��-lD����������{������ �-�@�`nD}O�\�)Hb�[P�FUE��9�v$��c@��/1:\c^��M=T�=�P'�ⶎn)F��.���C5��!p��yZ��dN�n�j6���C��%�Y�6��S=����ٞ�w���QjA����Jm�&��9$EW$�3��ث$���G�p� �!˪�j��<+I�%�q�qn�@��c��q(��w�N�7T�a���G?[tǝR���1G���q�~@�"UL�9QG��-�&�5A��v���]��CV�TR�.��3u-):�T����Fز���:��寬�P(~��{ 㤦��U$�{�8_7[xI�q�b�	8g���j d-�Q�o�v���8d�F7�h1S{�;'�iǤ����?�E��$���X*�@ݦ���Ӥ#��Ad�#��N�S��k�7d!�`�^]��F�����J�i��D0��[���N����X�� k�0�5ŗ*g�a�5C�m=.���� �3�]�m�U�����P6�
:���Y{oR�R��.&v���m��ohdV��S�J��з*9��Y��{��G� �p�mB]�|Yd�*o�5��ԑ��_�4oܿ�� R

Y�A�h�-�}���F���#J�>e0S;?&I��G�e.�*0� �J��c���e�Mֺ]N31`�Ʋ~�Ӄ��=XlxVHYEB    5b11    1480SH!C�C�Za��W���������%h}�Y�o�8�����QX]�2Q�-*��AYi�H�(W��N��g;NN��<���#����x'1�ڎtfB~���c��[�e5Bǟ���T�U��ȱ?�}z��PWO�f���]��O�����E�d��&���y#��LY��d���M']�fp9�GfY��&����Je|�o`<V��]m6��MeL@�H:�	)w	y��R���5�H�Z}�Cxl~Y�W3�k���)O��L%��a����Ɣe�F�|
z�.�<��4pҋ?���� �z��ٙq-`�����@ p�u���r=���[)��)�oNS�$�oB7�dt��kzSE���'�+�&~��=U�ԍ�r��Z"��u���7�V��݌���;�Sx�>��uށ�y���܏.w�?�6��D��TW�@B�4���2L?��ڑ�]D} ���w���E�܅T\���Y�E����(����3{�0Iz�R�N
� ��'�԰W5S�]w� �N"=J29��T,DT<U�!�@$c1��-4�6"+-�̖���k��SlC�"X���ύ��C,�����Z����-����=��e�<,�:�+����7Hfq[�����S(_��_aB�m�)�{���	_�0}w���h�Wl�1 ��i�[�-�����;�A������Ue�H��%/��]����C�0��Իsd4�����,����恆�.�К��R3Q����X���*OP^l-w�U�a��5B���1���t�<-[�	����%=?���D���U ܟ&f�6�S�b?*�ؤ��r��F.��ƃ�O����tSp���@c��=g��ki�z�x2P�e��@��S!N��gk k�Ҕ�/`����*�,��Ks$R\��C���j�`4�0R6���4vĪ��%�-��u0ӽ��-��*���t]GEqPB��y�F��M ����n8�`�e��}G�^����8㢿��m�L��Nz`Mt���pt[�G��u�<��rD�ίYl�l�n��NU:�q��]�z@�$�EoF좲�O9�d�:��P���Z7�?_��b�B�yď}�A���:��p�'xk뽴[R6��k&��W�t9�C�$-2	g��ZUYi��v�2̭��g�A�TE��G�H@�~*
��Ju�A@!4$�����Z��B*'Ygw}2�ͼ�����؅x�$O�W6K�*�t'�[,� �'��(�s��T�qsN���B�wj�j}��ظPU4DE�X,����n�Rۙ�{�5g�䕽6Fq>�CS ��A�4C��@jQ�+�.�CR��Xj�u��M�z���P�\R�0 2��;O_S��Pa���G/O�w1�	����� �9	����j�N�%#��/�;0������^�h9��]��b�p���m�(IಃTK�1t��$��c0����1+�������R�wJ��<.V�Qg��5l�&vP�j5����m�D�ۭsN���aRR�jV�7r�H���O�&W��U,��k�0�+��Z}�`�
5[��#��H��LЪ�K��H
��[��A�լ&�AXQaY��a�����u"�	����}�*�)ܰL�Ҭ]��zn�t	��Q1)�s��Ԙ������/���}'&2��i;��b��Mj���� p�.��3�op/��(��j�`O��V���R�z�U��Z�N�x�Y��ɈO��f�?Uਈ$O��QozZ�=����_�vG��{�S��0[��pB�R�Y�S��J�-�%Cܻok�uE�H,��A��k9�u< ���j�.,�|�����7�}�a[Y�ٕ�����6,�?І�r6����͘�u�b��n�ѭ�+v!\�Y[��X`��?��l�wvYF�s�bV��� �y,'ׁ��*{$;��1�����+W�N���F��V�aWH�51�����,�9o)���-W�a�[�V�͸2b�W��oϾ�̊K�2���w�;Xw���6$:3?���!��X�[M��.g�f#<>[1z ����J��W��M�� �k�����HQi$9(D/�@6�o�g3N����h�Y�u�����IR�������������x��=�R%�h��J�w ��L�UT�o�>�˟Y)�k�#�b��2�b� p�E�呛ml���Y��K�0��UZ/�j��S'�R���H;)~�8t�L(OM47��n @����E,p��t�ʅ��%k�Kq4��ݨWGip�>�98������">gKAC�߭zu�(�ȁ1N$$��F����RL:xéAV���ZҎa��ͻ1�0q�2Ev�n4�ru��Ch�g��<߱��$N�j״�e���S�\vB>Y�ʌ�+�l�DV��D���<������b�1�T�٥6D�٨aś�F1h��ؼ�g��Ce�SӲ�r���%�L�X��k����H+�ҁN.� [I�!:�yڮ���&ҕ�%dR�&;�b�h���pԜ�\%�_�xꆁ5�����4�*0��s��h/# ) I�vj>��e�������'Ɂ̚މ�c�U63/��&V��b9�v�!E�v�]u&e�PZ=��Љ��d̀�/=ce:��3�$��QnJd��Q;�J�(�7U�qYd��3��ii�02;���������D�����F"�I�_�-��g~j�����Vg��Kݓ�}܃����; �
¸��a�V�#I�OV^r;e��4������Iv�UQ�q�	����gdk�X�]L�P�.g3��d�2�I�Dm�}���K�ؚ;ϫ̲�K�C�l�%}�t��S�J8�a3�Ӗ�vI\���P�c=@������6��8C�YTO�
I���1/pX k}��/��f�7�*�1�l}��[�����S��=Mf#�8�H�͠�|.g�	�W���D�l�cs����5w���Q�5�4/�؏�v������`�Y�FTBg�Zs��|�f�������/�q3)�
��B��V�G��÷�cr	Յ����6�~������.2���&�$�Bo�F�|�� �Q�Aa�����d��6#����`_2�<�[�K���1+m�J�K�;ک�|��e��\` T�,���)��*�b����})��lԲ�J�OY�t��ϬO�~\t[Aɨ�����.�)�����Hq[G(w�/8�Cհ���6]Зq1���vo�3���%��➮$�'1��'c��9�ت"���uT�`�H��l�
R��Y7"8�� �[o���pwYfCwd��~�ʄ�}�ڹ��JȒs�0�����f�4\�Ƀ���\��EB������@OR���!��^��L+�"H�����~	E��˪�s@�����LK�2�e��צ������\&���fL	� ǰX�[��JB��s5��c��T�Q�d���ۙ@����k�F3�uL.R�DT.o�I�6��hm��z�۴~�i����3�\1RI�y��t�Y~����c-ɟCQ&��X	'��:�'~���������JYpk^��H�(m��sP��(�q4#�c� a��E�1ɫ��J�)܇���j(Q�^�FF��%:F�3�*��^3������s��fS�~8&I������sm��N��:�o�N�^\$E�~�jþ%"�
� 4ɻ#wF�?h���Lc��A�4��):gh�-\Z����}6"-S���ʧ3vp� ��B��Yٜ�˩eB; �p�d۶�+�� ��I�Z���I$�q�:��
����ǔ��:�f���y�]ʒU�.�/k`5_��u�]ˉs)�v�\�!�|�ل-d$����p[s�^���Ԭ�k�M��� �	�")�@#�!%��d[ꭃg��t�=��I��zjM��Dמͭ��v�ꇞ�
u�2F��OZqQ��r^^��跊 a�,�{M*��I����g|�X�p����!@��a�����r?�WB=*����ǽ�����O��y�6pԿ2�#��N$�\V٘�y��A� ��o�P�����Uz�<IA���1@БX.���m�PZ�
rDvm�_�^�<%Z��jc�*���I3��.���t��k���F҃5�/�	vFz��3����?���2��`��
�x��_W��W�J��a@��+Rk�I�í��n�[xՀ����`/��<����E�?��J���Z_������p�(H9�Q*`�dJR�����0r�j�������XH�E0�W��mӤ���`��$ջ�O��K#E���3VT:��h���=�ގ�q�K��u_��a'��HT"��+ײ�TC~�	�v�F#�(g���m�b�O��BBF�E�>�i��q�C�h;�!��,x5��)W�a��q���?bx��4"��W�������<o3���W��5�����,���l1+����9��
{Q���s��yj+�ݳ��,��&�M�}8e#)^F��'��������7O���]���k��t.J����d��S�Ѱ-'�XKrr��0��wil+�"D�-<�B|,���<r)oJK�����!\.����Nj�}�K�V�X�I���T���˔O�Y��X�>�[@����k$.�S���Й�t����b>8f�|2�f���{���ML�$�^�L&ǎ�U�.�_b���fn���m���wg�asu/�>&�`C�� �1�f�&[KvY5�E�,H6�ɍ$�BU�8�@�P��'ܐ�Z�M��[ը$��Q�.��ĸS�VC��_EҐ�X���H�WOlH��%�D����(��9�l���D?`U����+d`AO��S����΃��x��n��5�
�[��j5��/���^c�z��-U���vPB��s��7�����贈]m<�j��w�Bl�@�I�O�DSD�>�yW�������d�h���AA�k�l>���Ԋ�N���QXr���K��?��/������S����X,x���,�vz���+�.R,/�;.@�I� ,����c��r$f��u�a�kJ9;�<����=����5�w��-��/�`M8��䋤@�q�y�~���Bsq�խt����x��� L�٢3�ϺH�J��\�C��!�g���Z�^���O�M��BRO]��<��p4�[؎�
��`���s�a��#�2�[� l
�Ax��