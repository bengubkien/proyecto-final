XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����q<bx�ݠ[��ᆨ^i?�%�PuF��*�f��=��qȃ�xr�nf!:�A��.��z�лbm����E럙VA�i��N ���{��#�{���k��!G[�S N�9$Cs쏃yi	����l�$Y_��PX��ƻL��J�>����tO�?;�	����9K��SIɋ-���X �N�?o �v,�O(۠k����$r�㦩�h
ȍ�T������E�7�W3j�`Aj����m�I�i��%�CA5D
��@�\с�r������q�5�zWs�ZX���6�#��G��5�a^&��(�u��R����{��8�|�ʮ�Mv��?�~���F�dM��M[����Gnm��K�s����l���Jw���p�}3��؏b�aO閹�p�pQ3O���.��cDi�^w�p4ðPRƑ��v3�����0O#���;�κ�%#�l��l�|���_��F]���+iL0��>�9P�rM@=���E������Y�\z��g�"�������8 ����
�U�Z���D��-͙:�#��J�M6$l)�Ӓ��;Px�|���6	\I���y���&kK���m5[HJ-�/���U�ɲ�U�z�b!.�ueY�6�E���!T���^�d�߲q>V���M�K0��x!	$��/��K��$1��,�� hN��EȯL��ޣN}�E30=hB�SX�nIPPL�%���⁜N�nc�Vx`Dg�(�_&��כ��ZXlxVHYEB    fa00    31b0: G�z�`�^��O�C����ku+vgз��G�'=���A�-�xķ�-����������i�'ZXlh��!���Z����3�t�@��� ƿ���p�VaQ<�J����1���h5\9ù[g�C��x�`��4�x"N�*<�ٔ��}kN��dB$Y.���� ��	c�}�gf@f�Fg��Z4�����->��!��%V� z����?����H����pu���>Uf���S\͵���L
�sN�9X����W@��tu�z)��w��j}��<5#NA��WU�M���ĵ�áݱ8�Oc���-_��؄���Rf�������R�hل�:y��A����1���f��_e��"�]����c�� �]⨼�ff<�.����G�<�-�-�Y��v�u��]^2��h������*������9s��p�R�	r���5�.�2I>�Iӏ�u��p�[ E��ӹ��,�w��V����-?�(m̾c��|�����e$������{��[�L��	�G>W�����2������t��G}�6�O�s�dK�P�����LA�>!;殞�l4nI�n�]|�7�x�U0�n+Ĉ �~�Á����0[dQ�@]쉼sloXb�l`��=!w�]a�_�V&�	���7�[C߈߸�pU����>�{���%����}�-����� �T�0�+f�n��%�R	U�R!]+KVe�o���:�}P_I�'+��_�1�c`|�Ik$�U{_ƽ�\��kֵ鼏��d�w΢춴Cq���!�:2���w��-���A��A�P�=.��;k�'�Q����s�,�p��x���2��P��~���s�\��+��_�\	F�.�=&Oa�7z�Z]�CH.珹D�l��rً�7[sf�\T�����|�ī����O�Q2.���8�h�y�!X,(��h����w�;�S���O�4R]�E��M�:8>i%=�����e�%4��Ǎ�m��&]r�/�;�8?�	�9:)F��hf�B�A8!��b����^j��i��+��v�>đ�rN2���ӽD�Mҕ���SK)`*m�w̕g��^)�}�y:ѲUU;�9�z�d�-m�4��XƤ׎���߮t�T��ᘺ��oP������6�Uo�S슏�G� �#e��H1���J�Ր<w��CD0�^*��_TH��B�cA@�ۋ8��n��p���&)4n�����d��ݠP���6j_M����U�g�@��Q���(}k�4H����lO�,Ȣ�Y�՞������$	3q��H��1X";��N�$Ի1\�����$���z��չ}��?�F�l��{2!�_�������{�=U	b
!�5�[�n�)2��d҉��1�Kgx��4a���9�b	-\����G?$X�R<\Q�c9�s��%�D�z�`�bh����Hv����l�k1o�⚗w��PR_�d��Q���Xu!�U�i�K�K���EKY�v��A�`�|��:�5��g�u���Ѳ�NW�̛�\Ƃ�F�4�������P}'��c��r&�w�|Q.*kuq�`&N�ޯ��|�c��if�u<Y�j�-�b��	���{�a�(l(Z���P�e� ;�!���zQ�
��T�f���'��q��Hj;�8^/��"�7������CbNc�a��5�0P�uN��؎�k�ivl�,��Q5.���TC�P�[sOw"諆�z$���@�\��xj�_�y���F����h�4=�lSy�P�Y�F*��p���4I�/]E�ˍ�����o��ud�� ���y��i�}:���jP�u�P���R$��j��.�o�M+!l5pYm|@�8 t�TDg���(o97���H86�v�P�7}rH!�����l{z����i.%:�-����/`�sKS�o���D u��-�z��8���o��!�`��l�ׅ(��G#�-����Cm��0xBH\�F��
����[]������U�I�f0�͊2�k��Ki�d_{�Iۼ�d=����wN5B+LV{�fՆ�Qjo��
o�؈j�C����4 ��e0"��NkI���ۣ+Ē� ����іW��j@�w�J�Pc,:�*�a���V]MTu�Yp!N#�פ��pbPn���������;�>�쾼R5e�
��f���hX���l,�B�x�;ʍ�����w�}]������Aal�	#�Ɗ���{���$x�τ�	Ji�ֵ��:;�P��?�V�P�4x��b'���\<w�����VJ���k�c&=��	D^���uGI=��:Kz��W������F�� �u1'�^<G5~����*��`ς��X�?T0-[ 6֩�RJ�ʕm���Δ4 	+�-5�[�
��]L�PgGJ�n{Z I�5DBp	��_.�%F֡�cE%u�f�v�
���[���tl���ˀ�,;K�}�h8��=�v��!��<֞�{�|�{iM-ֈ-�w��3���!�����PĈ��oh���M�6�S�^�e�}�*�$����T[���<�L�dC�{\ &nr�.�g��G	o���9}����h)aTh�0�����3��\|[��������D�@G�n/"��lOҦ+1��"�9�@Ü=M��j5��5i�)�wHi)��k$b W8wJ]Ea���p��{�W.�����NnBifU�!��ݬ�Dٚ��qY���&,MR6m�Η�s(ʗ>�1��2+Xȧ���WO�+E$	D�j�&�YO�c�v�k��<��i��$8��n#�tF�`^l�(��#�[N����	��>��4N�/
3��4����-4��K{����/�YK�K`���
�������p�U�O�l��hd0��6��ª�fZ����+PxUDi�?�z#,�P:3�o"��2�Oc��\$+�J�F1� �w'���]H�\���=�t�bQ��d=j@bO?=�\��@���fO����(�� ���G�e�U? o���-�.z���h�q�]Ŏ���?��-������]��bA�õs
�k�Xk p_	S���F&?�, �uD ,��5�'��ےλ@M�g����^Ё9�o�v��u-L��B���/�M���:3h#��>�1�k�Ly{���E�:����%�����U��:���p������dP\ ��yJ+�!K��L�DH,��u~�O�[�ϛ#YDP:�YZ��z�PG���j��S�qs�+����-�̼���g���, a'<�߿�S�Qj��q��B���igVLM�*T�r^<s:���� Pa��B�B��z���z�〢��F����2w^�<_�N�֑ZC�Q��h�\���~[\?)y��PD�1X�K`���5�ُ�����W�Y�ӄ�ޚ�!/��ea~/Bj㓨��c�a�Neͭ7rg3Q�/�؇a��z��\+U��^�Cϱp������%"��܊g�z���S�)Q���⼙.-0T������ABR-ǀ�������J���y�&wr��1D�`��0�;�i�j.i�����H]D���H&PŬ�l�������y���]���_r����N��}h�g�)ʵ }��ƃh0�]��!�#�+�u���m��<�M���~»E�kp���ތ?ЮS��L��	.�n�ݓ�sW&.��50h���nD=��b���4m �4�9�u,�w�E/D�%8*�"�km�[L��QV��n��Eݷ��ж�gŖ���P����M�D��,�!���yO\��If�s�V|)!s��y|���g�d��e�Q>��o^�[h!�:Ǆ��{�?���o1�Ft ڽmJb%�!�k�nA�弢���E�~@�_No4�{L��~}�i���[ �}ّ-��AeM\̿�+e����c����Xun|��X�!:=y#	�փL���7�yd� �k9���ݤJ�	�Zͭ�z5�����@ka��8�V���-�Z��r�{>K�y�*��F�O�J�p�G ]�Z5��q:!?�����V�Ժ� ���gX��ꩢ��Kc[?a��;�$N\�T ��"��[������C�Y�k��
1�.m�?6��X�.JX���^�}�Y������g����1˃��\����c�w�A��W��`�aj��wtsrf y��a���naB2�no[���v��q��&�{F�>�mDO쑘����+�)�"�+	x�|����e��U��@JP�Ǫ�#�b�$���:��I\�������(��6޲�D^Xj�7T"�u=t�m�n2�<xZܻ�}�����o�D+���F�%�,�}d01 /�N�'��x������j �қ�]H(�U�[�a�#�Ť/h��#^��-��(��Cm[����D�����8ɔ����Y�[�}@�D�"��E �'�O�L�e���Y�$�O�A�����_;��S�h6�%�a0vZ8�U�b6�}���a�ڭE�|0�(��z��P�-�M���K�d8o��yj�x� �����!�ht]ո����G����t��ȸ���4���G�������QkoE�J�ɍ�)��r�]�]�@���p�w��?󂷙w/��f�����S�g-�^[�U������hī����Ga�	7��q��ߖ�f#����:d��<���fs���H��s33�5J�K��a�p���g��?�4����r$vE2�l�:�r�ݸ�Z]xaI�nr�/��
.lrq�B��#���~��p[��� &]�񺼰�����T0��]3f��Q�$�d:T,��/ vB�\��h�hc��e4k7���e�,�f��A��ΰ����^g�@(|.lW���3�=yJ����ǹl�FXQ�V�T�p��Wh����P�&�V�o�݆&�]��K�r��
K�jTuO�Yl2DI�1v��پR�Z��0Q�%�S��Z�H���nY�.����	b���3�$GZ|�W[�<F���lb��z�s��[Y�`�OP�S�C�g�<3#8�jN�/+�ݣg����T�cdt�i:�)�)��?6m���fdC�i��Xn��蝱�����ƹxʲ���D��c��o����m��I���
T���ɩ�Х�oC��mAA��yP�v�\ܠ&A��#�[���š�vU�h{C#��pY�2��IťaG;~��hB_�����kP=ˤP\��Ŭ��އ���C���3����Xv�1��H�,���%vh�i*_N,(����q�VIҁ��\�\�%�OJCN)pf���7Q7e��S�L��wjFy�9b����bv���jU�������7B�0��û<xͱ��^ٗ��m��8��K)e!ϭW-�3�U궳��򒧾ڿ���F��7�3g��P�N�R\�r�^�ePuK/9���9�k�̗��nw{'����_���gd
����߾�N���]s>{����;�P6�	��-	��]\�Akظi�]���]�)~��)�¤aS��fU��L�Nn�7eۆ�S'{�ʲ4�ù7X錝�x���6�i�s����@N�YS3��G���r��|~o�|\C�c�.Kd�T4[����}��TQx����4��opm��<�*a�Ə-�2�Eظ!}b\��ǈ�on6ː�R�a�E���\/���T�֜�s,$F"��#s�7hw�$�8�~�%t0�gx�G�}�'a�۰˴���B�΍{�$U�yΒ��*V! �vJw?ؐ�����\�v>l8���tE�
i�g� ��GqQ���(�S͏q��_,����ϼ�����i��7�ta��˸�j��Gn��Ȭ����d6������:�wU�,Y��L"�3�c�*�H�0Ż�"�^/��y�l�����3}�K����el���ob���9�!|*�B ?Q����!�-a��'Ch Tq�!Ī~O�%��=�	��t�T�T[���,r 	�n�"�E�rr*>�>o��=����� L���4D��S��S�T[15t�ƢT�~���V�u����`�-���x�#�0��=Р�'��r�S>]��OuA؇���*��&��y�8ņ]c���� E�����/^V
���B=������pV4( y.���1M�+~L����җ_�����O�mbH(l7ԕ���Yl���kP%�O��ʴg�>�)>Q�R�w����(\ᦘ���D]�G�^Yʝ�ڜկdR�����B�U��32ֿ�o8����B�����F��%��؇(�E�+���Eg(�NWے\4Iǩv�#��4�T����*�+D����ْ��Fs�W	QgV��hT=]~*���`��չ{
=0<)�M�͜��J�u����.���?�,�F�|ʰ�>�'
0&�l�R���t��2NQ$��}�`2C8xW�s�8����"�S��U%SĘ�<���f������Z��W}�g��=ͺ�����in[^<w�
C��4��<��A���塎�����ϓf�{��_��G\�3��`�]E�T�Q'��	-�^(ss�&�R���g��+�@L�a7G�s;��&u6��pą�)�]9�u�1�B��:�jO��DS�H�Ȝ�Kڔ+�8���Fp���� Do�!vT���ӡ2c���ڭ��&�)��\	��֩����rU�uR�cl�**��0�fK*"�S���x	�T�AY]헽���A��|���"��L_��Qd8l&�/��m4w-U"����W���y#�'ϒ���oL%����V7#_�A�6G��3��\e�4!�O�F.S{%�#a�����9��M�Pm�)�Ӿ�L�<i�]���gG��C��W%;���5�$�=����n�U����\�v�Uw@#��h�w�)�����MR�J��5e��~~5끋�U��o�C7��8K���y���%�q���2�Ӈ�ԃ훲�/S+7?����7ȝ;/D-��������#5�;�8�u4��3��
S
��j���l,M�����XU��ʚ0?����p��,LҌ/L �k��F���8���}�@-�0����,0Ağ�;8G��Z���溴B�Y)�����d5/X�B(��O��3$9�y,J�y�$cW�g\�6����f>T�m����3|U�)��ض��Wk^g��:૦y�m�F6ܓ����9[�{�l��y�c�'��:�v�V�~E�ݛxr�dr�H�ۦ)_@�a'RďǍ���l�?aGh�t�w�tG�`y�L�}�tl(����ٳ���9sҖNj��&{��0�;u��-?��BD뷜������5h��OEw�5��O��X�<U�}�������fb����G!��r�4��]?2W�L���Y*���zӯ�p�4�O�~���>G�Y/;�&�-��g��L��W廓�-(�2L�Azd�z�������@��O�L1_j
�myM��WO�Yܑ�g�瀥�+~��nF(��"�j�Z� 1W٣�mE��u��̼�R|�	����.�A
��6X����I���m�#sӳ.s�=*��`֝�̜y�@F�8W?��{�>��N���;��A�v)�J�M$����Eԓƥ�"�&4�,�;`��Ϧ�Q��y�ꤳ����:��d9�%�@�2�('�0aMUl;�uWC�+����*1ic�#�z.G����3]���C�,��áPN���ӆ��wt^:p>,�n���n	�Ž��5�H�j�5@Q呌���I7w5��vT��ƚַ��uZ� b	:��}ά��b�;�lv@1�{�Z����ck�><��{��I�5��W�Hڕק��)�f@��Sg��˅���H�W��E������D���I;�"��2I�o6@���W��8�F�S2��K����&8�IV��W��)c����<�Ŭ3��V��6���bם��G>�t���O��5�|M�}S]�1tQ�A�OV��R���d�v��XIVHk/��	�[L,����5���(�J�b>�s�@x�!#o���un����ξ�E�	�ڄ58H���-m��k��O[w�iyo]�Fή"��sL�0��	��a>s�q/0"�U����~�rNV('i��TJ���P���|i��gp���R~��w�p���_��<<%�g�@ w��tD6�;h֓���oH�sݺ���oNՌ��g��+��˅��v�	�\��0n�P��Β�d2��O��h�O^�%���(f�#(����d�	���3��*XoFbd�@�����M����O�_/�~s�a����.�f[5lo_`�<>Ƅ��XOC�P|R�K�#���K]�k�Y�� @1�6�/>g2�/�d�����[���u���J�\s��~�����тY���AQW�[�+"H����RY�s+�YP�������z��s�K���ʘ�C&ĬDH9����A܃��\�]iվΌfw��kmp'Vе��H�P��ӕWV*�(�ߞ�T�R���i�Zb��pR7\E�����lx���^d�ӹ8D���t ����>��J�e ��j:ѣ�`�\�dg(���W��ԣ
�i0��?iK\��|���B5 �9x�<��D��0T���E47gQ���=.�g�����mLn~|L{q(�ɷx��[N7�(��J�r�J��(��#�;��3l mz��zA��}�w�˿��"��?fU7�˲��7JOz�7�b���u�;O|��[X�����uj�ī��s2����Q�p��2����[M@3���G�B�5�@�%��p���&?���D|�ĮLKj��:�ϖ���h��W}>�޴���ڭ_b	F&/�}*kD��B@��HX�e��˔�����$�d0&5.�`1���A�Rj6Muq�![�&R
��+�pM)`�G�TG���ߤO'o>bi�h���7��>R��KRFn=B��6�Yt�:N!�M"={��q�_۩���&$ª�JZ�s�~>�ug�{�&8�:ޟ9�t=M?��ЃK�FC��Zxи���t{������`{�X?-,'XC�<�6�A�`�r���m@���1����Fk�e�A��\�@�s,������#�I���';���JN1�njr�n��#��q����鞎���%A���Z�]N^� σ�/̋^�[���T<�w�/%^miMh<r���,���A�kn� ��BL�0��P��]�ew'���ğ��N����C��$%��;R?�e-(W� K[v��P&A��>�qu����&��!�H��k�J'��>y��gg�\O�!�l�Rp��s��I#��T�q�v�x�\���i$@:�Ѓ��Z�XC�n
�-�#�w���n�F�QB�Z@~�F�qc�~����/6��M��f�����|^ ��� �-M{���<��x��h�=qq�zm��bO����]��{rA��GL�y�d�עK�=5�Q��:�e������̈��q���}���|m���~�ٞ���M�PZ>�%�=�.ߗ<�G�5_�&��*�e��ٮn
�m����ʭl^����tM��SN(����Q�M����#�F�m�Ve�G��͞� s���<�^�1�&A����������j���#G �SEk�bJ�su<�_J������ z�h��E����@M�72$�8�j������o�Mu0�L�Y���xy���^{]���!�H����g�+����B�6*�1ӱ*V�-��-�"�i�}�0o4ڡG
/���2,�m���O��#)ǖ`
8��v�2ׯ�@�K�f�^�*�y|���!o9�. �����b��i�D�钃wt�PH95<Y���(+�RR
��*g6{ĢW�}���F?o��a�Yˤ�;��0"H#�!�vK7`8W�yz�c���P��#�z�]�NX-��P:CR��E���;:�9�O&������=YX���T�4w��r:t�c�Ď�� p.�B��?u��T^�&�\��Vz"��K2y����2Y��ȂO��(��[�㋗Z��c��i�h�|�n^ur�S�ҪX�iz䉭��lxU����w����3�?����y���ycfR�!�1��u]La�uZ�إ�v��f�wI�$�������a�*���n�|��"����.�(�a�����~�L#H��:�-����R�������:�[�l��Y������{��ܩ\
m�|#�/�ܾ��U)�x���
��V�M�=�����)׆�o��&��G�~P�M���w��T��0M$@۰M��+�y�2�ɂ�#�.��)���b���� ���c�F$���{�X�P3ٓ��W~�!Dt�![����A_����b��,�6(�1 U8���z24�u*�h�[/��o �#�� �<{��\x��^νa��y��-���vIl�Z��=��7w����B~�s���G�����*�\����;����	���l��/���X~r�^}cvL)PNwdh���$�4w�Ww#/��J�K�]�&�l}KΨ��%�~�̎�?�^��+N�PB+�C"7q	C�����E����ir��#��`�<;��>�/��k�V�C ��QJ�39��Z(�d�q�܋�xX��[O�ߚk��D..2r*-BS��Ϻ�]�C�7vۉ�%����:��x��\���n�m�;��^��5�(�����|��c'|�����*�Ȯ�UuE&���%��_7�P�5���h2��s=�zD��rW���X�S�	���Ӟ4�v,'I9sC܃z��9�9�2��W�~M��o$AUc��f��q�ы���96k�ֲ�����;��%T��C�OΨ%X��{�*��D9>���9CY�.��<e39��ICR��q�U�Y?9l��+�hwR����Y澔��y٦C$q���tc�YEZ�pʯF�k;v`�����yi�� �]$�u�W����?������]<�BP_�8�_R�R.;_���{T�)$�)�۴�Q�}�`����528XH������=RQ�}������I��g��գ�HF����jL>���
�g!�Mh��1 ����5��?||���,�o�i�Y/s�L���yH��/��E�BX/��Ԅ��F��~V�@�~�s�Lp�5�Ep|���&'��֢ &�#,]��T���p�@g[�b�[Y�i���kǜ~���Rvٍ!��ƣk��#v�w����N��EhE����M�;*(�P�C��?w�55��a%p��G��:Ĺ�3���x��憥T��4����oZ⠨'JP��b[_��^,	@"�+3�fnAK��K���4���K|�I�Vsv.��`%�� @N�b�z5�0�{�(L�{��$�~�,;�vEs�>��\���Y@��֖S?�leR���	� sV��dbz�3�\�t�&c��D��)@����t�9ίh2��**Ղ�#�i7�"�`H=`lsU Q E�$_�4ڷ���V{�ʙAn:B.�U"��x��1�Z�$ߢ'=��4��̍�'B�B���AR1jՖ\R������E�9������bs(���S���V��R�`z��`޺��L�2Q1+����Y�u��G���X���C�G+!	��v���۳v��@��$��)�m�P���G�oC�;߄��[��ު��$.��)��C{ά5���bK�kp��b����G.Df���eo����0�_A�لx����Rv�8I��E���^�jc`	�r�U΃�O)|�3Z縁�f�=�����%��+��e[o&쁋�K�$��eŻ\j�z�\8F�"b��o���y��[	h���Xg7�Z<''�/g��]�`��r�Wxa���	�m��	��D&���i&���F���(�y�ilQ����� ^�_j�o�6��@1�֫S4f�ϸO=�@����ԍ� 3jy�gX��%�c��)�)
�5�޷���D�9��f�	5.zd��鼹 ��,� �� �	�a�㈤[���}'Q�:5c���C���>a�����"Q��]Ey|r0�c9�U�>!�`�X1k3�&p��_��M]M�l@�
B�=�1D�'�%%���/��u;��Ao����K��OzuMվY4�c��j�&�	=f�������I�Ŕ�G��\�l���� e����,&y�����o���;�V�kof��!��|���I��݆RN���PtP�����z:~=��I�%]#�\��4���F�1X�r{������]�H����j
� �7q�vD��)�FK`�ÔF;+�h~U"���dC2@��<�,y%��������*��k��j;7Y9�0�ܓ�O��	5�Ķ��35mOR�Oˤ3�I�1\lGP�o�ቦ4Ɓ僾��t��8ĝ��~w��Rd��($���0�귎A�A��������sY*����O!�ֽ\GT�B�8���lPR�9��g��xiI�I;7 k�{29����$�	�hO{p��K�O���<�4��֞kQ�þ�QsXY��þH������`��<��omC��pOrf��|�
�622����T7���Z��B]�E��>��qT��o�@�ڎ��������%<�&���hU��0�XlxVHYEB    18e3     640��"�`�vwt��q*fX ���d�!�?�A7�%1A��u�hY�V�U!a�|h[Us���'y�N8X�(�|	þ;��ꒂ������X5 ��s��˿hd�P�<SN��,�XmS˩4b���py�W<�4�CF-�s5&��Cn����).s�%2�T�"��&�[ 3�<�Q�����J��(�qeOF�5��
�[����$9D_��F�\�}�h�#׺6nB���������t�aƸ�������3?v�~�zD)C�-�V
ڡA�����VxHMd �>�F���m��F��=ՔjO��=\S��hS��3�ݩ���DkU,[��$������3��ߐ~�O�u�-FL�p���k�B���L�{���#%i�@����Z
�@[!���Yh��R���X��D4��ܵq�Nx��!�������~���\+���Ϡ�KRd�UC�Z zK��q���4�( ��+��C�<ުC�߯�2X��ܗ����L���~��e��H&��~:�T��0jƵ���.��P�\��q��W�����<V��H>t���M\�̪@k������ɍ�9�,V��e����(fC�����\r�Ҳ�~��ʲ�\��ꬴ��ը'�"r~U�P:���s���u�Ƒ5���1�é��epW�ΆĪC�wsհA�"��ORD�!u�Y���Z$*h�p�)�H�B�	M�m'�����%��!����O����Խ��z�0+���6.Xp9�o��������Xp��aA��1|*�t�"OI0g�g~��kD���SA&٩5z+����n���v�y����H�Ϭaq�X���q���O@�֣|�f_ƊE�>���9_�X䕢b�(Q\�];>G8aΉ[���Sڤ����&u_������C~��'�]6�Z}2dW�I՗�~�R���q� �9�9�ծJ�}e�b�>v�����Cr �^������Aғ�U�����*/~��U�vy��(e�|��jA���W��.=�_��CD��u�3�!0u�n�釢|w���\_D��#��}Q�q�6 qa".,`����U�;؜:�������o��r]���g�4N���t�y�7~T�J�Z%��MT�T��&���.l�1��L3{)=���������/���h�2��|����:QQ*�j�#����rcw�k�!��Obƙqi~�cn
9*�p�u��
�Qm�ل��/6he�-c�gQ� ��6h��)kk�g�On�T�bex$jM���8h>���(Jc�c��]$�2z,\�:��Y
m,4n��k�^���J�f)#ê�������^��E����ڎmBUu�����z8Y�����B�4�/3rr���S�[����RI�J�g
Pj�,6e*�X�~�}�5&R&���	�����@�M�l�&���RF,~`���Y�i�q2O|2Ac��\�!�x6��2�1*	e�/Ǯ������@�"�3�烇�z{�S8c�� .%�&5tZ*cs�$����m�)nu�\Tm{a\A�vB�j�	W,: � k�j��Ҵ�L�3�n���?�B�p`�