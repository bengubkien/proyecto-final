XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5P`A_�X)L9FoI�u�6k�$�M'q�v��W��m��g�Y��`�{�K�(����9���|�OV�g\C����p2'� x��i�~�a~�e�.I���܆�G	�a+1���Rc�@'�n��7��v���j"�d��hId���I���o~\��
�;�mxs<7f�,�����5���m\k����<��� Ցxf���i93��v�9�wI�LR��n�m�MާT:�B�@�eM�7����"����S�IR	�MXp�~��8&�V��ࣳ���ܚZH��a�w���]o���n�s1\�V7�}0�6%����,�h2���c�U8:����%��&G�RCx^eEsM���6HS�YI�q�{'�LL6�o����V�� uhғ�[�
&:��@/����� ���A�=�|�3�\k�աU�'�'�h)�7��7�LH;���^]g�g���>Ѿ��xAv��1��e��MvV=�����n��;��j���-oD|W�H;�,|_(��[e͚p��YQ�'V��4ç�� XN3�ԒQ2&���kto����k��g<�0��E���Zc\�Z�Ҟ�M\��������9O�� ����EѢ�Z]cG�-;C��jf�>4��WI���
� �'�$k75�,�j�H�����G���5bM���P�y�h^����|\�u(n��o�'��x�ׇ;Ƙ�2��X"�By;�4������L30Z?�W]TQ1��\V>F*{�E[s�/���8j-��.�S$XlxVHYEB    2870     c10�%=�o�ITZ�����m���h��ܥX�����D��D����.�R�q�����]J��G��D@�Vm��Z��_619���j�6����hF�;%�;x��3|�i>��z�}�Sj@����������v���:?�]a碾˧���+:¾� �si^��Q�����ڶ�v�\�m�Y_'������Od�]��H��������oM���E������ц�n����Kl �aR�B�����F�a�#��~�!N��j�y,�#H��G�]�;��L���� �C���:/z�Ջ�У��ut�[����T��V��7�8Py����/iX��<I|��ڕ��>�Ar.��:m��μW%��u�X���Jc�7I����'�eк��:�/oT�	�����'�(4�]�Uw�*������E�F������tNs?]���"�3�rӗ��zN�^�ow���b�{]�/��4j<�0���6�����O��[\�سc�n�)�o ����Mh�Wm��6���h	�}I��6�d8��X�E%���6�k���+�$��9�49�ߢM���A���I��l���!�FQ��1�Ԅ�<��alә�I���T�����N�n�m+�U2({H�̄�X9���:�{MV@�!g��5��/$��O�����d/0�+�)U���L��=M�IY=g	��� U��3�����=m��!�	���4� s�<;8�t|��y��Ӛ	�M�1����������̃*�{?J��oo����(<��D���TC���w�^��[��X�؁ȴ�-���tW�|2_��^�w����C�O�o!t�e,r��J:|&�FjkIq�ܭ oM�)�6����±�����;ι<Ǩ$��7	�MG|�~�LB'����Er�Ʉ�FG^���}/�=�D
���5�V$��=ĥ�3���f�yn�y�q�-4�D,Œ�oHF�ju�n6��Xrc����h~�F��0Xw��vs�P���W~��Z�Rϭt;'-�/l�0*�`�aZ�}�|�<�89�1j9O$����/v>�ݢ��e��F[���V�y�3�����^>����X&��}޹Д����$&$�)\%��
�=��mA��^���h�2�(R)M�<�{� ����6��؍�N�Pr^��ǁ�I��'J���>:,���4�؁33M���R}�HڌI��n���^a߀v���ǽ m�;}�F���~?�얙@\Bjt�U!�S5.�&�w��X7: '^�d�'E<�t~p�h��T��EfDS:0��^� ~_����ڰ�y7Ytp�q^�l��)_w&W��| y/$5�s��O�"���&����Pj��blέi�J"��R��i�3��ŋ�7e�X���\�+j����BE�]=['>�{�2z��9� �E���*O�����nL~��&W
	?��L��ʶXt"���sk,��cyL���ڧcB�62�/�/aK?`��<�{x�G?2 N1�"�|�q��(��y��2�m�=YBd��wb�ɯv1<�h��Y�B���ϔ
y��g5d���NGж*�]cg���qR��\�>Z����$*�OC�>6X٦Έ�� �@�כ������n�1c�s�ڀ5-BRg��#��a�5��B�Jz��-�g�h�,:��a�|�^qok���L���;��uW�|oz��c"���[ȧ�p�$�pa*>�Cp�Ӣ�c�n������+�1�$�D_n�حT�$��|DF��!|OI.ﮣ�/Aw�g� ��*���;�"X)�2���w�r"f��9|>�D*�+t�!��;����i P�3��2�h=��5�����H���lumLq�	�v��%�Њ��p�Hy��6�2*���7�yܙ��E��5'y���]�B�Qۊ�� �'x�>�f�#6WO���kr�n����#�@)�+�+k����F�Q�"��v�������L}����t�.�V���p]]�X��t���%w|p�¾����<<�^Y��ck�G�#�m��C|d?&9��"M��[���Ю@ԕs�c�'�-�FL��AO��Š�եS '�V7Fr��)�M�VzEƴ'	Ӻ��9��&�FV���_�i�)pj�Չ<���t�Px�\���8m
^j#�i��́�����4c���VR,���2�X��Z�ϱ�i����c���C:a��6��9~٫�G�&�Ҵ���ʴ�@YW|4��6�1��Ojf5-��|��_rZm��nu3��ݜJ��y�`��tʩpu �n�i��6�"�ж�I���kc�Ο9!c:e��n�:�TɹU�DwP깹�ے��'��c'�8�C�<r�~��*7�y�H��{��-Lh'�E�Dm�Ȏ���L)�ԝ�ϧ�W�:i�r�ՃzH���u�F6�r'c�,�'L�,��H�R��{8ƻټ�D��,�i��	��bP!�F�j���Px�����V�%�/Rtν:�@>�}=��E��X8�na�C+�ez�nC��Tm[7^�GN�"��;�o�
�"�wuRa�^r����t�������^�e^lx�#�\@V�,L��B�)�Ⱦ a�'�q-p��]����(����p�f���7t���f�t�[��o�b����,�ѫ�w�2��Y?z��� ��9hK2�Y��B�v�i;�I�Vx�43]?U>�F��[�G�6�[�2��<YC�6Ǿa܌rQ)��,�	�/����1��-nON����>U9�_`��K���z��6�G�>vՅ>�!��H�%�(���s����I95.�rW�g�׋�8���g��pL�Aݻ�
lL�o�y�2#������ϡ	�J�"ɥ���%!�]��&'9/��m�ō7̍&VǦ��M��rE�@�R� M-.���|I�|%V@N�K��m7�<E0���}&x�tkN���e�g�{�X/Z�B)ׅ#�>��g��c��� �G�/P�{�&����V̀�ۄ[ǟ�@(��L�H)� w ��Q�"��O7������v݊w�c^�