XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ۤ&*Ȱ�9�P�98�{r���R*�U����T��=�Lj����Ӳ�%C��￢���eD�v�i9S�z돱����� |]��b���]�/�#wgL�WT��ѡ|2ܵt��,�o��^2��؜�-2���n}���eٞ��n���Ƀ*H5��]8���ɤK��7�#�Z%t�dП�=�/�2]R������k���E����\bnӝ�����t�>��'vro��i�����x�ض�=X��P�����.M�4A��ie�ú탇s��S��5���钭+,�y�<m�Q��W�QֳtW�vo���ÏJ4�F��2�Ɵ��E�����뿐tV��>����Evz�M��h^�h�D"�Sϛ���m�*I�V�.���[�,�И�-7���}��]�Pp���4���I2'v�=��}��/T�*��O�(��7ypA�״��D����.�%�'Bu�X�a�OJ2��̭��X�*�E5�n������V"��[��W�)��d}\~�Tv:UrR��ߩ<j�lm�Y�}���+�	���z,%������Q_�p�G vCG5w��١�D}���k�W <Z��%�&t/+)���� �&�'Is���6{��6�@w�xph�Xm����N�('�y�mJ3ɑ�bt/B*r1�H],��nW�?��GpF4���P#bz<����}؍�Hw�T�s���{��H1
�l��Q���
� HY"���*�`�!�)8��x�\���J��6X*��ҐMY,�XlxVHYEB    1320     7c0X	�VU�W��U7��}�����u�fd���i�y�WJj�����aV�/Ҙ����dh��1�V��ڟ��	�g�R�i����"%�@ؿ�C��}Xh^���8�����ĥ����\s��R[��?��[���U�g=�cZiho��dh�B����# �u�/8^LOm:��V�+�û�v^� �/����`�-cڗ����TM��vH���~��r�.,
e"RZ���t��%�l�|A�F�4�G��(��1�k�8����������cJ�B��)hඌ�)����u��A�Y!��X`� d^,����bPc+3��"GN���Se�G��?��|*����`S��x0b��%s�k�d�Q��<�,Ū�rS�Yr3�*&�kg(�r�Yk<}f�s��v�a禥 �U?�{�o��v� �b="b�������zT�
�8�;�8��5+�{��s8_������G��4T����.@hxl�����;�$����	BNDS�Q�ųt�yag��N3����H�LQz#���+�Rzk2�r�aWyh�A�HD����}�Z���'��'�`�||RT˳=�q������dՋO\���3�7e��lR�����J�^��텂LH$bI!˖�	�S0�	R����R�RX�Z;b��q��S�w��!��rY��\���A���R�r�?�[j;E�n��,,2�γ
�<�K�RF��		6����D��N���N�;���*�s/8�
�l^ӂ���W�����m]�	� m�}wpF.���|I���}���v�Ѯ-�滿���u#�G"�Zp�ނäv����uM����ahh��������9�n��-Ƥ	�:Q��+,s���ҏB��� ڀ��Olf"��~*ʀ1����T���$�8ׂ�nd^M|=��7=��,T�#�f&��^��gs��v^(�/(�w����H]%�`�۹���Sq�����Os�� lzvVuK��Z��aT=�)"�M�dfq�h��.�f�k��)R�l�w�]$C�����1��)_����@?U���_�=D��V��U�Uq>�g<X��œf��o�*���"�&-�_�C�s�3jgc��q��|��U�xYD�h�����N�#p~w�Vy="�)q{g��Y'P��:�+R�M��ʄ�;3����V;^���g�m�'�9=��8�3��ɘ�R��ɻ���i���Ҳ�퍊�>z\�8>�ת?��bt�H�3kո��Q�¶X$0qx2�	w��#��{�Uv� Q��{(
��x2�q��C�Rm����*��Zڱ��� <��@wa��u=̂�S���b�Z�;	�E���0rC�]ܭ�6�3�[�,v+$U��<G�V,q�{�~\���O�P�9����Y�K\W�Wrz����J�����$؄��rX ���E�x������vj��g���� ,�`��`���dN7�5=���s����R�RЁ2����)��aWG��O+3R0��
�P=Q��D���]%)
ӕ|����@�m�j�V�{������OC�5
��rN�e/I��a��ɕ�i*d����Hj&�·�	КM8-M�9�ן�s����7>h]���Dc\s��;�gh�v�����cb�
��i�H�x:��aeћ�^��?^�|hG���Ns�����ɒ�*]o�\w'�'��Ԡ!d�sH�=�2RT��K>y�3zWv{����/�k������� Y��W�}�M�}$�D���xY�Ui��cH!�<���Ep3JbS�B%����2!\$T"���D�DӊFS0,3{��vdЃ�'P�b�ȹYVʹ�I	�-?���KH<���O����\�ߖ�E`��z�&��E���2�ǒ	�=q�m�M����K�z�Y���1GCp��p�0qx�d;�C��h��D������9Ҵ6].y�Cdl�թs����{ͺD]�v�-S7�a`