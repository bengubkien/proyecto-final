XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j��0���`"%J�Tگp�^��G�[
�Ǧ���Z�v*�E��- �hh�������sy}�N��P�u���♣=�g�ϳN¥�ӑ�{i1B�'�����ާ�m��K��\���̅��{M�K"��ƽ�;���Ҍ?
2�B��[ބ3c�O,D�04�ǌԘU�MJqK����Rt�^�u}Wܶ�9B�g���%)suc	7ӅE�ӜB����&Pq���L� 01����g5�|��~�0����M���zG��~AXq�4a�l3�i�m�o�u)���4�=+�6%U����0;��Β�������l�I,��t��9��?V2��tP�k��r]]GЕ�|L��9O��0�o�����'Ŀڏ. 5c����թ��+	 s���2_S�N}"u�����]���Y��l�+7���J�%��B��z�����u�恓?�)����ӖA�V@�z��x����;�a؈쥫W��(r��;; �'�`�A���� ��o�UC^Ԗv'=I������X��o��t6 �2�Ĩ7O���b��b��#���褀*�������TZ�2eq�9� a�Fw�EY}�	���";ޗLA��L�tK�o����4�k���^l5�<����x�7v��1(K˩����<���dn�NoV����
/�4+C
�L�Cr�cR���[��͞��c*p�IVX?$�K��A|}�t����6 !����@4�9 l�X)|	�����c�+��1���w�\@V���(�XlxVHYEB    61ec    1630�;��Zֲ�E[Lu�I��Q��ӑ�,<�Q��6��v���m��H"���G<Mr�TE7&KƄ�\�ɏ\�����E�R�м�	�VG|@yO�K����y�?�D�Ҩ�?�R�<A���U�����MX�K?p�@��.�j��]�C{@<ڝ�J�Н�f��-��Fvk����Q\�ѯ�hN�ں{ֈ2�w����bi�%o���-#�j�*ͯ-7>�qE�p	��&Wњ��Yvġ:+���i�����W�W��F8eF�Ki潳��X�ˏ��v@ Q�X��5���s�������	<a֤ǋ��;�2�����zq�,QC�i �q�u\+��ކѮvet�7��(�n9W��wc�Xe�!)�qj���o	�%p�s�,]��$��:�69���(��?�&;��'�	��;���#*Ϭ�B��
;}�M�P��j�Lx��<��k��n���%Y��I鷽,q	�@�a��J׬�Ş��4�=H��(k`��a LlU�	�Q��#��g�DO{�g�`S�1 ��t�}���l}W$j�F�m���<�*��穦�"� Er4�?�ԗ:Zm7�����1! 9�З�T
�_���G��b�wڀj���-�pM.M��{�H�������_B��.X㡻���Z�������4�S�|F�mH$���M��Q�.BAP�W�Uw��(Em� �%Q+]d���r��6o���D�;��c����N%G�EZ�6�}�T%L_u�䛹!��e��Ѡ͙�U"�Ё���F���G9q��s��׾-�Zأ_O�����iN^����i_"-��8о#��@h���-��� �O��'���8�
�k�����������ИK"5��ތ�2�6�"��AI��:Q�ˉ�nGxU�x��#�m@��]���0�w�	�{ς,��Ewj1"UB^�F�
�K�I]f%�CZ��-�z�ǚ�#�~n�-���$��ʍ_�،�#8e���.uQ|�#��a:a���2-��;�� 1�L�"}Ln�9���D~������䭼�:\(�.A�^W�Q*,�$�%�!"6L���.�f{�{����/UӾ��$,LKr��_AX���Aނ����/�!dt3X&u���X�Y�d�X�Y~�-�֩GG��,ݪ��H@���2ī��:+���_	��8�'їp����ݙt��l�$�Q���UQ���o��}����2���UҴ���2ݬ�����j�.�������5�ޅk�:����"�����~|o\Mv�2F�!fF�È�3�x����
�Vi04��/��e��Z�0��xz�?3��uE�^�:k�i7#���Ed�ĵϠ3�g]� ��<�/��HFvO����	t�G�f2�Ir��ؘ�s�jU%��铲��AL��3�\O�ͷs��@�ñ��`б�;!�N:��:1�=sls���|t�s��_s�[�-4!�@mK�Оc�ڶ�4�UHS��`�I��>u�K@�* z��4�|	�s���B��	~.�I��W�?�:������V�
��^��/SY�|�0c�����ǥ��E����f�����'��RK�8���8� L�+�J�c��H#��2�Xz�R���W����O������~E���?DM�hne��B��Tn��)��T��C B�E,O�j2��hx�[ݜuB�C�.~�)W��T6��b�	�o� O�������6
o��r+IJ�ł�@��+��Dz��YD�ԫ�ݕ �ٞ��a��A�F�|��B���`vV8�û)�������K�)�dF�j]�ۓ>N�E@��._=�~�]�OI�T,�)�ժl�̢xUX��q�#m��"|��j��fe����0��T.�����A��.	�4����I�x���e����I���
.����Y��u�W!0���t��/�����15.k��zHh�qn�g+�cvCe�3473s�5k`�)v����뀴	�:k"�c���t��*a������w~��o���֎�K?G�����~�o��z��g��ݴ}�ܵ>��o��Y�B��K	�i	#l�ԛ��_�\�wn>}j@ҌJ�9���T���_�b��m�o��(� �ː	DU;W�f}�AF��p`��:����#��E7�tmR$�,��6&�:ԇHI�@Y��� `�S 0��"x�v_��l�S�����/{�2Ґ�W����*#��W��������Us�sA	��KIJsݪ_��c�l��;�#�ij�k2� �nC.�/��}�{>�	��Y�a�������l�j�7�N]��|���}|v|�#��75�z�3�m2�`�'�YW��KO��'t7�{�O��S����@�Xz��#I��3�)W�����Yf����$T���T}��%��(Y��z�E\�U'��^�%�G�z0ft뗳YK��%�z�)k���7�ҕ�ND!�,�g0��k�b�q~��Li��a����o?5[?֒�������8&rb8�X�ʡ ���U��z���B��dQ0��u5~q;<�nt�XY���)9�+BnÍ�9��;TдG�M���\"9Mpֽ�Do�?��^x�(r��F��V�^P�m�it��8ʱ9KB�P������-���1�w�C����-}����� LnFӎ�o����uͣ­HATu�e���ĸ?W���z`��°;�A�Yp�棃�<Y��� M}�/�u{8j�����6���m=7*�M��=#��V�qtU��{A\+
雪&�Y����nm����z"FTt,�l����oe�U�"�S��,��F���s�.{��nV��!g�y�@r�1�8qA�'�����	_>
l�|�'䒄_����V�&8+j��k��8���k�̪���yMM\��&���Z�qW��t���/�b JQ3�B:�M���8�����fYqd�k2�X͓�+^��eڀ�p�˰��(�����Ĭ�����r����+O^��wn#b��(I,��X^��t5��R^�[ؠ�Aψ�gG�~T�r�_	�|"�P)y>�(�>�s����6E}�}�����T^���M�m�0��PH4~�#�����agob��#�&Ń����U����>�M�M���� �l��Z���ؠ�\��'�Zu�G&�5B�b����?#��@
��`~����bZ47�Q�t�g�1�� ,+����Y4��"S<큆�U�a��\�ө�� E��m�,j`A�w0��W�?�ENNt��������˘]�z��fe<Qov��9�w��r�io���<�b�`��7�@���I�����Mm�_�:�oD���W+ߦwt3ޒ�	��������m�r��n�SaG�=�*E$�N/��ΥGrY7|�U!/do0��`��شKX� �3�Ea���C���};9K������ ���t�R�M>nƨ�?���Z�cf��"��w�]Y6
e�FJ>hp�P���8�!�O����*���CC�=�F�ҿ�'=�Q��T1(����67��[�;��U���3����V��|;��U�]��4�ODԣ>���ά]��$<lA'	��9v�����O.F�'rf���������Kp5r1������<H�s����d[���}���i~�Ybw���3c����p?R�B�8�&��6csv��R׃K2�������]��L�qj��>\�C���mǃ~����~W+��;Z֬��v<�~�Jl��Z�D�������$���#�>`�QP-���3x�v6�������J�~�]���Z ��RR҈�Ytf��i���R�N�7�B�'���.�����BƆm�YB�Q�c�~�Es?�%{���7�/��*90D�K��+q޺�ƅ�1�*k=���`�n>��@Ѽ�6�O�S�-���:�@J&qw���=ِQOAv�\�m��r�7�i���- B)���|�����r����xoT���)S"v��:�|��g�d��=;iy޹w����g0e�^tU�0?&�N�0:d�'R�uh)�?"�S :��g(�l��iA��&��u��Y´Ԙ�,9 ֲ�K)�� 0{jEw�q�m�^�wzPN�gk-5XZDr�蔔�\��8艉!���=����s��z��#�̈́�:(����/��Q;��4���Wu�a�bv����H�<��&�V#��{u��9���J��f	�bO���8>'�W���}=��"Tҟ}��
�2�<_�ur��Z�Lp��t�B��Z�4�����Pv�w��i��o�:dd�8���,�=K
�L�qO���^\#����$MH֙"�:�� ��4Eh*L(v�\�`K�����!q[�h�VѡD�0�$Am���h��<i��-���Ǚgh;����%<��T.�s�1a���e�8�����9]P?���/~D��8�|w�l"H���_�bt�H���9���e�ՕTu  ���G�ܰV�f�6����n�G,��+�V�����Hj��ob~�z�`���T4����D_����d�*�}*ܗUܹ�^>�gc+�v$8�:�D #/�!�����C�9<
�_�ËharWx@k�C�-����<JNRo�:0�"�l��y��U�/�9+���G6��(���bh�{f��Fl'�Ǹ�����Ώ#CV27���<B�F�'�n�.VGӤNZq'}Kdi��j�I�;0�p^d�!��#���W��>z�㫤V�\D�6i�K\f+��FSBsd�zl�H�w��^C��J[�����H��ci^��_B�@/4R��#ٳ(�a;�r챷����Q>ĸ����������p�7'��l��x�q=�v�by�f�M��h||.�η�ݕ�:lp7cS3����2B�Z}O4�P�`���L)��2Pƽ8�'��50~J?���E � I�M{��������M��3�I�?�]�!�	C#�2Ȋ�`D~U46�$I��l X��yw��.q�c���l\b�A�jO��(<|�x���\��1g�U�~�^U������ؐ�3]�C��!�"��I�ª�3� �)bm�R�0���T*2��11��'�Y�����B�\��>u9&��/s$�)#�u� �3*�~S��������a,�	�=ӛ���A�y0��y,�M	�6��߸��Y(�N��D�m#̌�>E��k��'�pI:�L��!po�_�m�������(z��s�M�9�y�$�n}8��;�p�{���8��92��3���Q �c���mx��x�9�*��n��Kt�l�;ᅲ
��t34\���p�,\ڪzw.�����S,�`5v}��39�:��W��Y�B�p<����E]��8ΑdF6��ٟ������\/�����!���x\����K&s���LH,ě��_棧W�S2�T%���hu�;�\l垳'�u"�.䛀i�E�ٰa�ב���B����t��Ji�眽��_oO��"a�&��隿�!>�{^q-�w�N?��O��t��p�g��-u��{?`�r~�2uP�M�6V���1�[�"%Y�>�4�|�yH�het{C�Ť��nB�$z���X�NKb�В����A0��E