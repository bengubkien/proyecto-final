XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A�ְ% ֧�Me�Ue�d[΃�9\��܊�P�Tx�'�9��N�.�d����h���u̸�3��
�'��\ �f"-��j�W����a޳083�Tw�B3~r7�A��N0�����U��*�w��_8q*����2b���@Ϗ�g��$#@ߟ���$�{9�rܐ�>Ώx�Om��ҽn�F�;nνKl� ���7�A���;"��V���W/>z��D��ZI�{Ө!�tHQ���3U�����2�# �`�&�����=�/7?�Z�3
�|�u��A>�r�.�� ^��=�������\w��%#�D�����ճ̥�5#}�������ʍ;�܈zB�k�Ş�4����V���G��{TЫ�[��2O��Z\Ȁ�B���o����@D�q��1���t�n�(���@��T�kJ��D��]\�Ms�$���(�갨���B�m�ɼ�wv/�ާ�����aL���Q�i��.�#��I�7?�C��"W�HΘ\��W��[%"��3��/.�29yr�N'�
l#��nY�>��t%������AG��|̝�(w8�s:S؋�&�~{�r�K�ǈ�������PKُy���S0P�4|%r�1��El3+�~Cl�7wd�}a��.��0������f:e�W� �h��h��D.�n�/����p��V�%H��y�T5����
Bd��8��`o�/9�0Cp}�V�\���s�P �5M޺8�6Z�9�*,���Q]_��[��[,�SȚ���XlxVHYEB    11b3     7c0��w���ij7���v�T�J�>P���~e��܅�ӯлg���OC���A��S�;i��%O�GG���Ήbш2Vf~mu�9�}3��Gܒ��tV��iOA�3#��R0�3�n[�{�Q����"%�"P�)J�h���$��C;��5F��Pe��-z�������(��� ��O��9����fk�O���&��mzYe�������
F�\?s6��zOP�ؓ��8�_����TC%PI����+?������E��N�g�N���a!M �!��7�3��es�p^�a�"=����S�[G؅��	��6,y4	ǓlW�b\����a���q
Po;��"�a~��<"yA���>�S�Uk�d��|�����qo7��T�Un��-%���5� P��fC�i��]XT=p!�5��(#���F��(�v�<DM䩑�p�o<l8�i�97�RYω���`�{�����߄�\x�;�Q���:/C+�W����h�ct~RA�Bu�t�A��?��1̣B����pq�����K�-�*�lp	����?���{�
��w@���\4�64!��T4W'7�hx5j���p�oQ� %��(-O%��XA�ZpN�\��a���[�ӿ��4l?(�ʣ|G~5�j
@]��U���?`2��kH���R��@�Bw��,�F�i��7�y_��4�J76.���t�w� �'+RGnи�-��ЌZkq�ۯ����.ʿ<�lc*��@����sb�:3|�����k�L�>��'�t�3���"y���6���s_��3�t���[}�S��>s*ւ���7!3���Z3kR�P-��@�Ҁ ��rt��?q^�8U�4v���i�jɛ��t8�5z>fi�`7::by��l"��ܨ)5��,K=/O�� �O�	r����EO7���W؞�+kE5&�HleGe�ТfS�x����pR2�Oaxe�Y�`Q¥}�\X�[�?M�)֦�鵉{���o7\���l.�|G	�1Z4�I��+�0���X!w@�\���OO��-9�4o��w<��L�dP������:������DnO�7�O�o}̶��ov�q�/�č<i�0������ʙ�Y�����b5]��8��/idq��TS�fɃJ�g"N\�?s#�|f�V�r�S�+$����U��s=<D��ޡP��c�z�į�7`�Yg]~B&�k��t�F~�&��3��������z3NbcIs�ܼ� V
*l��|QV��_P�7j����z�
n���T Ф~��5��s�a�g�㵛�	�	����2S�y�("0����OyԒOcP�}�����ub��<����c��q��� j����8�T����5%�+J~D8mD�B����&��G�&�P�LKS��#wYA^�:�,�ո����(�l�*���h�c(%�luT��N���Q	/dku���T�������P�'�|��`�E����!�g���z"d`�xS�}��VbA%12�$Y���(Y(	�b(�$k�k�)|I��8)a�p��V�s�ć�����$R�y�1�*yǭ�v�ї�?qȮ.�l\��zV��u�$����+kZVH�g�w
�0�[�%�9�zj�K�&Z�T,��y��8�~p��iY0+L�����g��l�R���`��BI�G�S�Ȏqe�]�+Qjq�`�h3'9}�LA�9�B�ͺ�kX�Dd��.���W8��x�:[�1փ��������id/sg�l+��I�ADD%MY��.a��V�����}LP�x%�Yu�z7���b�T��=?ۀ^҅�Q?Os%�8(����b��L��Q��������z��͕U��f��iǽ�I��w5�B5���(SsIwfZ�e�(m~{	L��8XP��9.��C� s��y.~	���g��&��I��m8�
}��g'QCr��>	U'�U�f��Nǻi����O���