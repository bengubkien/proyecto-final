XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i���9�{>����������7�9�s�����å#n�1��Jt�����^ԫ��K����"�"�+PH��x�Q�s��1ZLx}��Q��X�� c�)�R�z��p�EC��?����V["K��ĵ�׾6�������{S�gR�]��VP|��n^�o
Y9��ሤ����z�� E��ṽ1�xE����gzo��C����U<�S�ݪ�n-��?����m	�b���ҜeG�	�Z�gTx� �C���%��=�ϻ���Z��1t{-Ǔ*	��>n ohF|{�0���.��,�;�N�AxG��~�]o n�R�(���զ5�X�>�;`&E,���<�����E�v`$��{@c)��DCE�~�^��_JS���N(�WX���
�z�_U/��X�.>L����%	�=�׺˯���ջ&}#�&W��B��~�R=:�����������������7>]�sv�v�C�,s@��0�ș]��Q��_���`��<CV��G�M�hF\_�dI��ƨ�ʨ}�'���5,��_	�nv����x�#�|����+�ܥ�J2K/ѽm�H���M��֋�Ѝ
kv'x�22��]�1��~lR����Ď��E��Q(8���Ӭ��7�GD!|/�sw��ZV4�����G�-n$�J�ۭ}��1VDT��^�o��e�W�:� ՅJJ���6����h��T���"X�['���X ���naL�d+M���*0��(Ɂ2J��Z�zr҄XlxVHYEB    24a7     b90��I��l}��j�/x򔳬�s~1ȞbI��$S� ���ˁ�7�Y����4����mr׻x<�Ɩ9���ixGmK�f#��V��?�h}�
�X�i?��]�Zm��G%k2W��������re��{7&�Uf�S($ o ȫڨQ^W���O9�(��jX5�."��e�n&��S�H��]t�A\[M����5^!k���=�s�2\����X���p�!(�"C��<�쟦]�����R�V7l�
�)E1.�
�k����_|�[;Ρ�v��/ڄ�\�+�7�
����c9kB㈼�Ek�\�R�,��YNv����&����;�������ƾ'9�I�I�-����|�C��8��"p�����Z�Q�/`m�V��f����kD�D�#��l�2��y�M�f��$^K��?+UTk�6��J�r��Zv��rO"l�v��A�{T%�C���V\�|F,6����xf�ڹx��oV��I���R=LL���<=l@��js�1�i��a�]f�B��2���{�tK_r%cO�ִ������eU�2�e��k����μ��X�=0�^ڢ<�)k�y�"�xG����]��"�
���t�Yp��ػ�j�A�"^"֮0�qj�L���/-0�j#���N�=�G�޻}ϓ��_$�K�?d���*�T�'�*e�D��)��{�p�h�]�1 ���aȲ>��}��w=�X�XS���?�ܚ_�ℒD��y���NݒZh\�(j~�@�bU�A	����G��t7�P(�N�3�����|ֈ���o�VسD���?�q�QD���㛭��m6�PJw�N^w2q�/��>B�zN���T>j�9��.�&꼭1�s�h��׀��K�?	ʂp	f�|��E*���:�E��s^gf�$f�0e�`D��U�����N��R4ġ�9������E2C��I��>��|��p"w5L)�f����6�ݶq$�s��bf4���6 ˲��\|�V��\6�SPقln����>Uݻ���?��{�3��՝v�5}����<� v��'�I��dNH$N2��9!�L��d�C�����~�j��y��mL����:e0,6�o��v�.�sjO�|؀-N�����OkE�]g(Q�덣I�0���T�?�˯2���n+�����<���|_}X��H���\�<_��V�K��su|�6P�#�hA�}�W$�������FL��9Riϸ���G���磽V�5gY���g}G>���C."�[�����)�}�RN��s����K�x�X����.Z*S�<W�i��n�N������"�;�~��e�Wn'�n�/+S~;�zw�av�7E�P?;J�*?T`�JXK5E�l�nݤ��	��������z_��;�8�1����o�0�(Ӏ���S�]߫� �u��cL�gZ��XI��C~��0?P�Y��6.MD`��3`l�ȷzJ XY`�W�wH���2+1��i0��������6<N���1/.���g��k����3{/ug��)�H�7ś˾5��s��!�do/W��rT�-Y=}P#b+d�I��9]@;C��ݣT��{�6�D$	h �fx�r>���F��y
����Rd�C�}��UCL��[O�˻Hq���I�\��c��vm=���녧G-��^�"���� �{�Β�B���r�������23xo��T��Yd'���1�d#|K�>X90Bc]{c��e��g��Ck>8lzA�x!a ����h��r��cZ|���y����x8���<����D��i[�<��&�WE��ړ^^d����ϊ"�.^�������ޗ�C�n�Ź�����iH�d�kU:7I&sI�Q^e20�,�ң�ॶ5tB�!L�#�ƕ�P�q�� �{ƹ�Fw��*��[j��2�E&JPaۈd?�"��ԫ���Ϧw�"�����,H(�pz����s��?���Z�O(y�tÖ�R=��u�l�f�j�5��wSW�A�A2`Qz-5�KI2*~�����NxI%E?`�3H�f��q���D�*鍈�������2�˫�6�-I4��s)o�'�wJ��;���1������p�'x��E�=��Ң���D/�=zT܊<J��ĂD!���9�m�O�]E�%SS�s�����)'~��B�Z*�?��O�Vtߞ�Kq�*�ѦL�l�`k�9~8Ϥ��w�Xl���VP�^�9����]�1����"�Aï�[���?����}U��V	Nc�¯��uA*��\�6,}�\�vI���` U����WVrvO��o+�/�R�ӣߕҤ;O�w<�|KfC��Js�-�������f����gKR��� 2�B{~�<����6u�$$m�a��_�p����'nu&AF�p;̇
r��ņ�����g�"�`%��!�߫��F���̆�-�񉺐��Y"�F�)US������s�n�:������f�6!��5��'Ǜ4���K#����
��>�r���8ť�~VOF�z;����ju�{,%N�����| P{ӮҞ�2�h����>��������QD�"(����k&7*1���{^ng�b�!��عF�U�p\] E�5��d����R]�,��Q��Q�� 	����i������g�Wa#MA���{E��㮵� W���fP :�岚9M6�e6����oux"���.#���Ma�u%	��x�)l�4���vR)�<���(и�N�Ƿ ��t=�ӆ7��務�|�Ű�IQ�EM�"z[�t�#�!4͡�}��	��i�hMJ ��u߲�aP�q�m-��*c��e0�	�u�jЛ=[�8R��c�Vmj�����C��h��_�xjtvN{�\�n1�t��Oٹ^�ObbVm�M�83��3�p-�:�<pK�3