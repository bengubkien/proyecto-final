XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7D��^�e�a��=|�'�IJ��dvm��q"�Q��I_!�<���͢hZ�m���Ce}�_	΄n��']xx�p�E�w��t�C��ܝ���B�� ��q�ί���)�ü567�{5�C]�͈O����d���'��T��)SE܎x'���޻=�1O�?��Ju\w%�,�2��A���U�gE:�?=�U��a�ڐ�;=r��A��1��R� I�J٘Fq�ɛ��n���{F��F�ZB�� FO���`o���Pa���sH<C���[���B�YV����-ʙ�$7�L|dz6z�M�6`h��}�F�_B��k����W��C�����:�	�\�{7^P�{E�w��B~B�7��\��Bk������E��ؠ�uus�����ޑ���]��X�>
���R��>q���T�q�Ԍ��5I�Ճۍ�W�B;�s��@���_��U���Բ��Iiļh�7��M�H�;YYr�+\����X����LOt�@��NˋmF݀�Q�uc[�y�����d�ч�T�H��&ͬ�8��d�-cL�Y��Cx�ݢ�jtcR��_c�}J�"��J���1�t]�F�4>y!��;�����n�"��Ο�J��H���y�z-xWu�2�Cᶂ�0ϥ|=�UsY
#`�A���>��,n�W�I�O2U��������|k 4�#I��O�B���E(P�7T������4�D���ЏOЬ(�q���Iڙ�~��*��h�XlxVHYEB    902f    18e0_\��t��kIe�0���m�R�'/�j��Ѥ��I�J4t�'�RHmc�Z�3\����ՆXL�#$h�<vR�T���{�U�%>�Ÿ���{hM&�����%Y#�����%���gДZ�i��~�*��XˮEÏ#0*MU�K���R�-��R�&��%��q8����9����_}#���A�pߦ:B�~��`P#[���#�+�PܷP����>���9�����;�ZL�:E�r�;IJ{�x�|z:������򓡣)R�f���M6f�~7�U�&?{$;����$E���l�xw���l�\[".�1�&+I��ɂ�zϬo�S��z2��ܙ�r��l�^Y��&m��nt�>�<���ʥ�hZ��^�=�X����{$��(U�p#���+��4�$�Z6��%�;U���<�7R�?�����7��˿��6�1����[Q"�`&k�
nCFĢ*�l�=\���)[�'�\���Nukc�Bc�@��j�#��9zK3��U:��pShl�{�	f�*�S� �ӧ��vJ����j[hX�$��}8�<�~e�p�5`[�-�%B��X
@�˂mDf�ƈ��6)�^���Nޞ�i�.�!�Q��D�ku�V=�� c���}ȱ����?�����O�3G~�S�ĭ��PΊ�N�	vΎ=�W�nVS[C%[�Q<՘�}�l���Fy^5��f���Qn�v�FH|[�/��%;0G�ñ����5� mFzU[�XU�8T�w`]��)�c��w��qB���t���,9��;�R9�Pl,��|�U*_�����);�C�K31,C?�Ӵ�S蹦z|�E��t���B�-bJ��yH�q8���?�c���;"�H^v������(N%K��ϒ���4���e�d"�mD=X��D��*�t��#~���ii���\ft	�^k0��!X5+/��������r�۠��Ҡf�F��b�T���H?K[S���Zɡ����4cq��4мU.0V&f�G�M^>iI�\�hMi���p P$�Vw:��J��WE�Q���km��&pb�BB{�J;���]r��u����pF�;�4����;k��K%��C�4�d2%�z���\���3���+Bx�t\g$�.�;��!	@T3HHp��:����|�st�+x�K���p�Q��c�#�G������ g���y>2�.�U��\1oyA�^�j��(�g�%rg3��Y�~7~����:��R<��Ùۇ�~��!�OV eX�1�X�%0s�3$�NT�p��8��x _�i�+�ƾ��������[�c�:0�\W,'��`�đM_QLMcۍ�B��7��ƀ�t�!)��t˸Æ�,z��pR���^�N�] ��q��~��d�Ɗޑ�E9�
����?�D?�%�S�m,�W�aX�u�D �(U�ˮ%��%�P���zK����0w����l�;'c�6��C3�� �.�e7�7���7��[��6�'\>A��dwYU1uaCi��~j�$�ڶ<������9�ظ03�K7�
�C��s��:��&5��Ǚ5V�,(&����B!�>�.ǻ��av5a��~�o��H���B�5Q�f>��R������[�/��{dv�>�l�W�p�{���PSH�6�9_1������o��ȱ�2��r'���W[d�X���U[��Z����#9%?��FM�(9�7ߌ$�[�[��I�Pޭ���Ic��O�:jV��:S2��o��2��.�*�ei�u!�hh�yA��+l"� �]*���y²@���M�����&A4(�B�轨�	��p�m��P��rO�A%�
����r%�g��34�A�w%\�Q�1:���͙�/���f��COm��W�c1*�5 a;��	:u��͙ʸi ˭��n#j}�y~=�җSU0�ʂLGg��c%�܅E�g׻i����<"xv�W����PS�3��e�$�w��|g����^�Ӡ�3g�g���P�&R��&E�܋KOIbLSy��D�ꘌ�s#mO�4sn���~ <V�@m9�h[?���z�.��cK�i�;�7Q� ��0f��M��ی���i��"P�ጩ�@��]�A�|���̰��32zfrL}�C�v��� �\����)RP� ��kh��]u/��3!�3���|A�������y3A*�w�U#l�ʓ��im��Zp'|oE ��E����O�8�FUG��<$!��`ɖ�V&���(�-�F`���	%��wuct� �ln�f�5��g���>9��+�:R�X�����^��\zM6K�!� �<�2]S�6'��|H�"5%-���qS�0��Ck���Ǉ]��N��#e�=�R�*�����6i��"<��O���f��&r��+��W#gi�xMܳ�2v��9:��l%]{�����Y]�c.VX�@Ajs���c�!Өv��1��� A��j7�%��nJ������#srA�=5k~_fԛ(�������z�wDY��������u��pP�;�w�0 ����g��}G�PC�*m`X\h���X�Le
�p���Q�v������h4�^�����%='1��6�jaS�SeR��9�1�D�8�S��jN,������bJyM���-!xkv/%.�T3���.ZФ����8���'�1�pP�1î�,��V��m���3�J���K�����hbױ�X,[���u/���H��י�}�e���=�'����!��eEG �2gW���(�l�DϴFtedQy�DNΔVT�u�Y������ (���J�B���d)���w��P'�q����j�6D�Q61�È�W��z�o�eZ�۪���Uz���������߄�߭@ٱCҰ��֗&'��T�8G�(l��z>N	-mYr�a�,1{�
��Y�~�X�`�!�P��.م��R�x����nt�A�	�G³�I=�
��r�d���-p��yf0]��t�i�T�g���NM���'.�[�GL����@M�QY�ǁ7
�׮�F�Ϝ��u���ܲ�-n 
j��ƑI�y�!ܮD��X�������B�u���G�U8�3a��Nͬ�O�e=�o�n���S�Tх�������{�}{���m����U�9���jN0l�C-�S���Ť7��8F�羖pb�hy0�8A�.+&�i�f��G]�j��O���_���z��(���uHi��� �"Ox����`�]ӊ(�X5�t��6�����o�x��,��q��K^]�:�އ,+��Ԥ�;����!Ax@q����c��G�^����w�6R���y�<���z��j���X�闠�p�ᵣ@$Z�����f�7�x�O�O� ��O�����5*
w3�����l�x�r��󆏗�z������gW��H�
�ʅ��[L.�D�p11-^q�<��VdHV
V����)6�9W�����B<o���?1E��{U�̱V^���+]����Mi��)��5��	�bUm���VB�d�a�|[PfW��9���:k_C��ts �����@P�[Za�����7o�RU����A�.X ^�ڢ�}�zS{+��()j�qaߢy�{��0��U�I��c>�I�x��e�r*q�P��`��E��7�=ďt#��u�y���$. .�G �F~��-�2��uLbUg~�u*���n1�Di]ݰ��_I�)���uq����Gb�XO���:(��~d��V�2�=����m��^�?�O�,����c,]��Vvr cǴd73k��0IT�U�C��r!��m��̌Z������h2h��=��s>��P����jM����*��B��&y��kN�ɫlKg�^�n��{���˓���y"L��J��zM�5��r6�6���aQ�Z�؜(Fn@����=*l`������XΛ�..q~���Tg��������$�o'�=A^����9�,C�U�`�-���MOۆM�(� �M�A�P���-_�)�)�2֯`�N�߳y�BV�iZ���]{y����6�񩙬��%\����Z�y�%.�ز�~����l<\�����?�/��>m�ڠLA����e��\�O$�?[L5�������h0�wOr�'pyi�B��{�&s�_A��<��G��^�n�n,\Gs�5R�+t��T@kT�:Br�XۨT��ogۆro<�u��uMF�r�=�����U���bg���i�
yw"\B�E��X6��"���|�P�iqM�\�mU�J�!�e:w�75��z��頄��D��?�=��09�gCit�,Ur*S�K��aE�5<aG�^cD#k|��f�+��D3\���ػ���$}����L��yr�~%��W�#a�: &4
�g'�m\�Fvv������4؛�5������,��g���礨vH����/��`aQ�"7O�Y���dc�;��)��vV�Gؕ�����4�Ё���򰢝ֆ��*���]bЃ��,:���Mg�ʏ�G\��C�P���~�P��� ���t�CBق8Ps+7���t׾�ĳ��r�PLj��:���.�Ru���ۥ��俭ѱN��C��������ͨ�LO������vAq��<�L�
������˒��?�xO�T�d�81��|f�o�*�r6�:e�o��׵�(~Ê�sxI@	�u�JJ��,2�s� =�);�IcX�j/�`/1����c>L[Hd�]2�ƕ�!K_��C$�ly~�G���G#�Q�;q$̇���+����w-L�ٚ< ϵX��=��׼�	�}9{~�'�)w��_|������i����*o��>����L��t_}Ljj���[�����[a%댯�m�g \EUL$+���(9�é�he볏�<�.y�Q�9bw���e��P��|Dt3���:�q6�PGU��	��G�d�K>���<K	<&�����i��>㤋�h�(9��G�#m�j�s�C]X��3���^"�az�S���|����)�Bb��1WOY�q��	�l�ZԀ�����h�ID������NS�OP _�'�f48����W�:�9?�D`TW��M�nC:��T �������#��S���M�c�����_Te�')3��f����d�5/�T��R���z�s���(;�
SdG�+�.}cX�ܫf�ct��h�W��R��-���e�-C���o����1fU��$m�'�Խ��6�W7I���UG�t�O͡�,P�@�$�*�_�Nl����qP�1�����j /�&N����W��4�=7�L�g�!,S�R/h�l�XK��<G�v�#�;�?y������E�����`b#�������������M	�>��1�k��X�:���"@��`�/y������)��8��	S1��hG�9���&�b@�O�NK�[��)�"@�� 6\����n�����<�̈́�,=fnt�'r���`N A��C�n�W�⃤��4:�˵+yg[:���]2d�M��j*�KU�J��sz��tc��k�^��T�����$�;�'�@���B�qE�ûCt���Z#����'2K���"ӗ*<t��u�ӳ�-�+ӄ���eH
������J�~*|�vL��	I�[^�\�Б^5�􃼛<�u*��?I���(QZ��;|@��]\��}>�n�3̅�ÛKPx.,Z;���E<�rd	Bd��uoG�4����K�UVۜ��lɹZ�{���)�#'�/�|�f	<,<������=��wV@ $��s���֍�,�Z�J��@v�}�»�7G0���N�2M��£?Ʊ�%"Ǘ�*��6B?l��:��,~�����+/��A��I"Z��	��BB�́T����V^�1ZdX�*�`̃�c�n�,��)K꣗�gg4<&�t1��������@�{�4�-�`Z��o�C��gٹ�[�LlʥMa=5�X˝�lb?���c�Y@b�<�E8�R��Yӵ�[���}7=�!}��3��L� z��F%�@��3���r�ge�cئl� {4���L�r�CL7�^�ʡ��<b�>0�jg~�4p�~���Aclz$x`��J�_K�P?��&�3�XOi��.���}ʌ� �Pl�#RL�c;n�'��2Kq��i��s�ذCUf�H��Z�>�i�9�w�8Y�S�)�� �Of(sΤg��W�R��o��� ��b��(?D�*_�΋h�ſ�#�a>�/K��>k��CaMJ�7q��B�q|h��2�'˕��RБj�q�j�