XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A��F�L�����Ϣb������{���}gf�{sӓ�3���=>D¹���O�ț�+X֙ɉ�@�_��T��������L~�,��8�ڸ�@r�7ǷǀiȌ�����)���R�58(�ٽe�K|<��Vn)�Z�[sKF���ȱ�2�9�D�=�p/�~R���v���J��\��p��v;��O�١]Ĉ̢��{»զ�
�ޔӴ����m��r@J�I�4_,��]�!Zms
����y�e�Ls���%&��nT�ȋ/��ʇP6�<��	�>&CI@�UQ3�/�/��|�u�8F.���U��3Ƣd�SL�.�o�F܁���z>��]��.�' ϩ�L�X4��S�B���Ҭ+�59U�I�n����L�Q�J] ��F�J�$R]�3a:r�YZ?�j�C,� �������G��Ҍ-�2Cb;�T�^U�x�iٯ��p��ڈ��E�Ѓ����{�.���;���ڋ�v��Z�W9�ƻ�|"#�&s��C�kv� g]o�C^��(�.��)�^��:i���藍_��ZW=�k<@zBB&�eѼSs���&*=���7N@��Q��n�7A87Աj	{�%��Ճ�W
2�D;}�,�t�n�l둕�$��#w���W-��VwS>\��b�WrP]m6Ň�Uc��� /Yյ�3�2�撪�����1�-3ì���ߦ� ��m�$����fdQ�ym<"K\ٿ�{.�<l�EY��Q�v���d���������g�\����XlxVHYEB    324c     ea0
x�uÇ-���@��QBӀ���!�~E��7�{��
�ʁݷ3��J�w�R�5�R=�<��ES�GS���Ɉ`AE������fn�$�2�!Pz+�yK�%zڠDkv��QE�cHk��$&�Y�*m#�=� �-��������Z��_[��5�!Zw)�����CݐGCs?o�Ċ����Y�J�"��iQ��<ij$��^��pۋ���}A��S�ItS��W��\�)�r�������J<+����{��F	hԌ[M+m^B�X�X�r��o���z���LӋ�����1%���
�%-hK�96���eCa��ͱ��Mw�W������t�m�EWx ?����\�5�ﹸ��p��~
������ݲ��o�e��ӻI}
]�T1� �p�ц�O5V�W}N���N��" Ѣ)xO�{���గ��?nbnr�]s�eS�T1�+�w=2�j�ۊG'�E�sڎJ�t{�sl�ۿKsdPdhZ�7��,&3 u��1���z���!�����}�#���x}NbySW B0pRf���$��H��е]��{:Vl��M�r�uLN e�S­��.��񰚫�A��x�sT���kU��}+L
��~7�����\���`߲���O�&�:4);���_��|�&��>���K�E�.��MYrl^ ���d4Ys�_���/Bc��.mZ����0��#�Y�`��R��v����L6;���V����ZG_�Ʀ��k�nu����B����ʩ�}�l��^4h��EE]~����1�y�$�b莽���0��Gl��O�;����.
na���9ʲ]��p�ӫ��!�V�@�|�e�*L�	��M-SCO/��Q�׌��I$a�W؏�ZQ;�)eq�^���_a6�����0����淒�o]V��t��QwCע��aT�MЏr��e�����V[s�9�Ղ�p����ͪ+�'��'�4~eOpɷ�f�^s��7<��.��3|:����� �^e����~$W���� Oȋv�[�AS�����q�~�İ���Êhc�Վ�+�+��UZDr:QS�G3Ꮕً#�A�@��<�5I����wn���0���kR�g���6�zS:�
b�g�;3GbgB'�S��ca���`9?i[��s���.z���
� �[R�K�Ȍ6��a�b��������y,7������K���I����@`N�X�Ζ�}���?Бő�w=���I���
�a���T��d���������E"� ƹ�{ܸ�����&�Щ�?�T��L��ŋ��]E ��{�D�l`?+�P��`@��xWT�=e�SW�C��o�v��|�GtSo��Y&��B�_��5̷�����XB��П��wk�M�N�@�a��<ĸ����A&���	k��=�B
���$����e��y��K�Ϸ��H�*N��-���w�1�b��*�F�g��-pc�$�l����&���-��Z��k�rԟ�dO�F?.$e�`�z��V%(]\��E��]��{_���fS�Fq_Mϋ��ո�� �!��~JG��KH��z��E�B�`+���''ȼ���N��q�d&��$����;F���ƲG),��=l��9S�Ip%"+���"�%�րX����R]�>I߂��f`$�,U~ �# m���=�z92!�UW� ���7�y�L���7�7d;_z�ͽ:P�����%�&^6����P~)ᨁt˅�JV��W%�G�RT��G��߸t!�(�b�o��B��`��+�)~ +<R�u��A��W��΍+K�Ϋ��޴�}]���m�Y��(x�Dz����g�w
�sx^h\��8)9�;�) =�L�p������h�9Q��ήG�(w�	N�{��*x!'t�%��/J�R�'�IDt[�T��ݨ����?��PdA[��_,�C꜎��v�۾���}Ad�jԊ��=[#�G����"��Z^R�R���B�o���<�3fG|YL2Q+)Z&L�B�e�H��W��SV���YǦ����jt�<G�d�d���̆��JK��/�� v��F���D���$��P����p�?xu�!���OIH���jVr�!�#:���P�l�\����2f���L�E-���:f�h A֙0$۠��R���?� c��R;�+]gDڞy������7�Hd�
���j�|B��������<�Pm����@q�1�tr��)N4$v���6鞰n	��T��K[~�ϐ�V�+z]%m-)�T* �_�O�	���5V@ka��"� ��W��2���-3��E�v�A�>��*�%�1���{�Qla1�K�D��Z�i������Hյ���7��29����T�
��z��,j<��m���N�ď +;D`"ڧ6/�����~rU��Ѯ�M�D9�@�J��������bm@V�or��"���S�|u�Kf9����
�Z���	���m�{�6f�2��~�,�E�]�p�|@��t6l�q�fn������U!�ꧪ#����IHQ�=G���l�gX�dLq�IB��᫐^��Am�W*�O�����
��'�vY�Z�њ'�r�Hd�v�I�#o�W
�{Uk�4B�@�$�9�5R�ֶ�� �˸3jg�d�{Ѿ_����b-`�O}�������r_.�%�'�X.N���:�����at��z�k68�%`Db�	��Hg�V�u�k@�u]���MP8�?]�OOrՀ�z(��UJ�$��#_�d��d�Z(
�ꌡt.��&S0|fq4)��k�>+;��r�.F$S>��	�be���dR�O�2&rr�T��d7������˪=�eb��-:c�gޥn	��)�
SK���z7�H�ݱ�j�0�i�@ͽ��S6M��oS	M��!!�U?�������y�O�g�v��N�߼�$5�7	��E���gt}���/��WB쭫��e��o��6�&Z���FUz7��T���5�T�Xn�X8�6�����><cW�=j%���RZ���/¤1�m���#��\�w�k@&��И��mx_�#���ũ�yN��1d��m�cͬ%r��m<�l.a	턯�7NL�xϴV�$(i�<��3�PO7	�so�J���-�v�'��̔�虧�
/2�����y4�b_���5��3QH��t ��/����~�K ��u7���\�K��{�2��l��1��&O܎YNyE�����D};�&#9Ós�ɱ�_b�F�m�8�ރ�����.����I�(u�b?3��k��|���8B1ia�_9U��c*#�����M�f�B'��9�v=��2ڟ��!;.v��(`,�F��Ҹ��J�{�W� H�\�u-�X�P��f��8��~���N����L�	[��\uePl(*����y����{n~[sY�K�4�� D��l���*�c��/�zY�h�X3M̊By'�ԩB(�Yi�������$��T��s�(��n58���N�i
n?ڶ��t��kgB�dj�˗.=&��w�	�c��&��V�k�
����]�Z	��Ƨn�3�o"��17��e\?H��&Je�~�i�� ��)�N���ܗե�L͊�~b+���9ڔ�ԝ�4�T���]!ō��$��D{�]u%(^�����WE@���.=���ί}�n�o}����Z