XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$�sC0`�qp�[n,5�>�P:gl�p�'XP %������WD��p��mW:T���׭g����w�R�Z�?n>,�8K��'��r�C^��ۗ�j4�J:�>����։���e�z*�C�qҥxHw_���x�zP�4��86+U����N5�X9��Du�����8�4�C��x�) �f��VC�㹁�t�{���FzfX-u�KC���*t�g��[�yfF���4}�,ir�K���4��9�a��[|���$CRu�7�p�� ET`V�]���J������B�-��w�
���ض��5jL�j$u)�AL����,�/t�M���#��[����Z�g��Y�=��q�z�C��`Xӄ��_�}��.�ڀ`��kc2:�9�?\7*��ܬ�{�����qC}k��Q% ��K�����;���Ie�VT�Q\�P�������@�y�9�K��)���$?�%���ͧQ�d���5�{A�S�O�}Tm�~�~��Qz�E��݃�ih�8I��N t�������w9tF�п��5���B�Gd���0� �B.g֐�A��M�h��x��1K���^����X�&�R�h��>���0~�%�^���g���]D�~��":��{v.˝�ή
k��e�Z@�_@O��f��|$�8�X"0KY�'Y�F�*�*�wE3�^���4��osm@���my�Y��%=��4�B �{,|�����9	��-��XlxVHYEB    a67a    2020����a�l�g�ց��_G�6��A!aUwq�o�����ya疤IB���J[!���(=�u�#��� �˪����0T��Ɓ�7�z�M*� �axv�7�J뫞���8��L,5��3��+'H�݅#pr��\P���2��xfe���F%\�U�p��<Ǫ��	�m]�}k�ZXI'����Zʱɮ�l��A@V�i藅�E�<	+�M���:L�ؓ2���Bl�hP(� �3�oCXu�q�1�N8�@\�[�ޟ�c�f����;��W��@����+8&�ɇF����JZm9u�Fh�Z��Z���3�c����q;��v�f����q��V�u}@7�,�\~������?s���8�X��2Q`� ���/�T6H��L=�w/��#�c}vU��q��wn��8��=Ml�qfx�E�����z���L�W�L���CP�=�o�$����QyF'a�/xRv�k�/Z�2#ĸ�%�.~�|�j��U4��!��>��}4�����yM}�� oB�&.����__D�g6�*$�ap>V�K��(�cdP+�B�&������4S@�yg]��p�����	̍B�T�m�E$�G�&���cJ��i�C��a�%oΫL{�a����Yf��LdxC�N�(��R����(F�מ��n��d���>��
�QH�Q1ǰп�e��W;��/���X�9��8�xO����M�����ܜ���.��팈���]�Y]��ح���P>��H�
�p�VR��,=�ir����A����sԲ}]�&@�&gW���A��Zf��:����[�� U���a�ŏ_>���lo �_/�sA����Zꅈm+܀/�+�!!����l�n?���||24��RnG� EH� ��N��@ȏi��x�]w��dTǉ�F$��������.�����)�*�ނ~]�� ڔ��w��7���ߘ�V�����.��:�.�?��A�7�8�v5$ �n�J�O$��H"_�_�B+t\��k���hv��@�k ��o�OD��g��ر�SP�K����*��X]-������^^.̈�ܠY�dO�K�*
[�����8{�iB���GR)��_l�jt8���$I�6J�K>Q�,G���~oh�z��>T����?�tp�����M�`�������GʘIO���(ͨ����p� e�(Hu�0�u��B�L�,�U���}69�Z�a,�Ř��;]�s�7��_�/a��%+|�-\�G^"�Q�}����!���u���a���}5+Ԍn�r��:L��N�[Q�BǏ4��������T_w����4Z?���E�\�K�|v/x)�N�!����K6��x���x$T�=l���,Y�V�n��~�ۜ�|vf��'��B��6{]���C�����m�a�6b��sdS�=����*���'-iJakS� ���P}
��%�����`�����H��_���F�����A�i��B���f�/C�������<�����0�b���t2��s�@�
*cڋ�N�ʾ��� �O��s�]O�cmz��~�)�:
�"Ҝj�=6�M]w�I��^�e�����Һ���{��晢ل�R������bm��.	��Pl���~��ſ-��J� ����ŬXՆ��r��X��ƾ����p"�V����mׁ_{��TH ����6�׭N}eMX�[ R���n����{e;}V܏k����p�����+]V������4�o����ܷ!�;	\?8�~p�(�U����3��R�L�`�ۜg	֍d\O�
���pp�qnK}�Əs�=bU$��z�˃^��4�^��i����[�뮄SK�=�^8inJ��:� � �k��y�&΋Q9�i�u1:'8B惵(�K�Y�Ð�}�50�f�2��iOZ	.O�=���QXm��N����.��%���?�8P��'�<��|�#����R���h��.���P��M����pX��u���[������=��P�F.�8�d�~�6���f�9(�ܘ�t��0,8�27l�~9�y�QZr�!�(�=NLF{V�9Ҷ�L�J)]{}�S��Z��{`M�S�U�tD��벥w�%���}�č�c�G�l�f�<��9LL���[�'h�ԲQ~�Z��F,!������e��5&����>_�蠥j�t&ѯl����%5,�X+̃�Y �͔�|�s& p�8�{Da���_Y�ntxNM�69�٤Z�Mx�����K��ܶ��e���I,
wǵ=��D������Ւ�r���DG�Q��T<Vi磍��Dk�K<b��h�1��=i9���l"UMLBڨ�t�������Y<_#�=3~�����T��.rױ�Q��炷�xh��A�Js�A��|�gZ>������<�}rp�bkl�	����5쯫��k����bT����A�/�����%�wW:(ce%��:�Rטd)�,��&�=�y:�� �?��v��H�/��H��jK^JI-@3��d��u%|ø-
#|��4֏O�"����ZJ��9B|���\=+�%[� ���t3��<3-u�W�-���8�$G� ��w�T#���DJg��$�~�w�Fz�~��W��E�cn�`ē��U~]�O)�V5����H��$��&��dF�QcT�B�Ś�]#=dB�X��ZW����+92¹���>�c%�a~J*"�B-����Aܲ�T�6$���Ui�F���wf����CF�~��KuF㑯���?v������ƤBv�{����x�c��?DK�fۅ��c�(����z��o�1'������2x�k�hS���W��>�m�+�Π��"�e�bkS:�mq�y,��Une�%�/��$��@�U�'<�ۣ-�.��m}B��3���N��D��𭩁��8�4�Ń���	-���R��x��u|�2����R�� �{��J��uv��
ťby�&#�aS/)zB����p?�G��XfN@&����()�w�\un9�Y_ӧeZ5��K�|����/6�Y"� �O����Ú<#jB-�6�g�x�G�O���3+��ۿ��.�?BG��p��+�/~X�C[�-O*��s�%���<���_ik8��Q¾R]��A�����~)��){q]!u��c�֗6wu�,�y��.]|���Ryַ�aQvv��8U9�"�7��x���ހ�^�����c���%�^��< )gwR+���E����D�_ۍ���M�GK~(>�#�i�k�K⥽��e�0���DcD��+r}����K�Ѽ
��Wa��ג)�_���eU�W(�:\}���P�l [�7%����J �Eo
z�>�0篢�Bs�'E��+}#󌶱�ĳ�V|`z����̫��(�m4�b�eX�[�)�f��H9�?w[�`�c�U��e�7qϺ�3҄��� ��؜T���PG��yٴ��Y�7�/{����'�[�FHA�����(�����%l�L��>;��k�Kjm'S����ۡ��
�%�ry�sK��K٭L*\��&�N���<�H�^�h��4=X�����H0��ڙ��M������5<���{S���a��"#�B�i+`g�Gy���_�	u�c��)�c���^	����P5��"�^�AF\n��!�Rp�_1�'O�9�?�9�qC7���*#$�ۥB�j�ݔͿ��F��$]2��K'\S��ӯ�n�}k�-w��Y\&W����t�_��a+�B�����N>%�[��J�����c�Bͫ��C<��[��ï�A߸��Xrf!/�����rmW�d��G�l:����	��C�X���@T��l���6�6��X�lg�����K{e�AHs�1{{�`��%���V`�%���LI�Z f|����9�c3F~��393���nk�/�R쉯��(��kgv�^�^��	(����ؑmѢ�i�\Sf!�-�e�I^��]X���K��[r�*�L����u��隕�w�J�{s��پ&��ȅ�D����+�{��Y�����!P�V�;�)��yR�6�P��x�ŭ뮲>}���dGT����s;�R!׳��W�f��L�8�av-?�B�~
I؉�j�p�O�"�R�ݪw]No�^4�я ��d�]1P��Dx0�	����ie�\����1޷�-d��'tsQ_l����-QYŬ$7L��ՠf)1|�!�-�l^�,W�c�My�n�YMb��-7q��.����X$���J�b37v_6)0�Y?�&w/lp8p�_�#k�r�A�ݻ��g��b��$��
�"�d�tt�  �!��uI��Y�3U.1�U �����_~����qWZ�:r�!#�ǏL���g�����.']n���J�Z��R�fu�Sm�T��=�c>�?�5�U.Y~
��(O��f����v���h��P_��������_Lne��>㼭{��g֤�zaƌ'��5rP�mx��,'��� ��ρ7E�M���	|Ovq]�N�"S�Q�*���<��_qLIQF4�~��-�>�]3���d;�A
�
��ԷN���`~~�0e���ԺF޻���ZdRx��܌z R��� $޳�^�m�~@��#���޻�h�"$1��g"L�+�*H�c���؈��C��>1�[*������iz��}c���k|�Qy�(ԩ<��
AY9h�Q��2�$�O>qӋ�fɌ�#�g3͋��aN5�
��FJg����CE.%�[�l2͑������Xf����ˋ0��:5Q�uQ!/� ?�K��ў.e���1��� t�v��B��fu�$�$%a2�ō���wr�N�֐i��~��#��sJ�7�ªg��ͩ�%�8�lWj�?!���;.

�������B��Ǎ�n%hj��z$�;��꜆�'�Wƶ��7Wv#�`P��=����#��4Y���̘o��ь͵��\��v�d�h'Eu��X��h�.P}]Tvê�P%���c(ډ\��\b�Z�c�1g���Ҏ4�E�OK���n��7V_��F�)�$eQ��.P֑������ �&����ή��.���{\L�U�S��-��H��yp���L�3��/C�*����f$�?��<��֦=���ڐ�<���y��/�ۘ���'=�q�z��O nUe[���:l;�P���_��j�-�n��j��MIZ�5sg��2�'2�Kc}t�4ajm'�3��L��1/S�&B��<�B5��n�4�tLl�c�i���Ȃ�4�	C4�H�Qq�c���wZ���I��_i(V��b�J{,��,�o�z��`n'5Q���_�,8[�Bu\}wNJLFꋽ�Zf'?U,g��h�(���:�X�*�^�;8ym8@F��z� {�:xT�o�=�e�U�}�{`��u�~i+��dI�?�h3��S>��v�=�;l��$ ]�j�
�{.��|��V��@췚�f�zsH���ԁij��^w ��ʋS��X����G�ꘊ�}"e	��1�\ 0-.�=��n֒�0I�oz �G�V��50N�I���&ᛜ^Ɲ��8+�u��5�q�C�fH��z�F?��a�����~G��t!� vBʏbae;R?dU����_O�0�ǢVQ}����S:G�=8��?S�cW�z�>���C|�G �{U�}ِ��H�OQ;��8<�р�ׂ�`xG�u�V5a����p��Ca�F�����NÐ�_X������@������I��rg�B��~�{%F�g�ts`l-����G�&�$��RL��kHߞM��,2c� j��6�xv~uSTR�V��jrY���²�psWx�;cV�x2;��FU�3H��b�6��&㎳t����آ�$,xs��(5��I�ʀi\AH%Q%+g����T��P�{�6eg�ͻ�0^��튏ǜ8�PۺL<_/�%�%r� R���}�Gh���/��~���4��g���~�X����ĭ���o�dH�[��X~w��+�'.A��A��^�D�h3�2P4y�FRu��>�X���E��7᧓D������*=�y>�Ng�yM�t��Ut"�D�|H7	w�o��6��N�Y\bR��]�e��ֻ\�e̿��=�k�'
G��)��x�1jJ{�bێO��|��u�Y�0���RI_��ޕ���PI�e L�w �T��؅��(7���~�����Q���)9� �C��V?{�f��9����[x���^�i����n/�$���rQ����H1�K%x5T�*W)�9IU�|m��Ӯy���CGY�OzEk��,�,�1NL:i��/�s���ݪPh�i��|���V��tP̰���2��6�L���|-i'�����W���y��%�b��i���rK �e���ƹ~��pyC y\�}y|�rk�j�Iri|�SuRvis�8SZ��gD�ˉ�Q�T�ϕf��&���{��r�-*�T )y�u���tL��C�S��Ա��g��xB3�ם���My�p�����9��<@tgD�V���	D5�$�\o��e�J�Խ+xS���K��H3cQM��g����q�P�J���`�����J���@��7T� G~�5�Q���� ��u���H_8��o�/w�J��m��͸΀��E�@䡘�Π�y�;8swn;�X���
�'��{���쬮�g�XɲJ��oG}�֗�*aݨʥà\u_V-�=Q�7ۉ��\���t�C�(�E4� g�8��X_q?9U�S &�0��P�h� �ݱ �U@��f������}ImP��/�'��<�w}��v`�h�����yC�jz8He{�>Y����*n��+e������[̈́�;�>� ���u�K�-E����V,�5�zN�]0��G_16^�@B���Y.P�{]�ڮg2�Ș��uF�K���ņ�����9D�b�K�.�׌)�-"m��l�t���b����oYpz4$�XnZ��%.��~?^uа3z�����;�:�ư��͘�����ި���z>O�X��P�[���D��p��|��T��%���&|�~L�K��m<3k�6$ �b[D�$�o��WX�,��?)��ĸ�Ej��g�P&��pP|��p�� �@��.|S�<;RW��r25\��(����Ȭ��r�7G���6P#��^�F���zI��Ar�s���̼Dq;��*�_���o�3���uxʀh��PK	.�_ac>�����f̓���e���K>���WhR�&Zyv��7DL3i��8Z�~�u���������'zPT6e^��	@)���"�N���);�I��:Rk%�������5���{xŴ���P��Dvv	�eZ%o�?7��on<�9���C5۾�Eff�x�KY�g9E�<c��.Dꔁ��'H���{IrbO��+�*��?'�	��k0�)#3�Hs*�l��P0�Y�2\oi��F>i�PO�Za@Qޥ�1u������|a�)���*k �Q-�'I@#������{�<�#y���t!�2� )�!���8�J��t",	���m�]�_�B ��cWO%@�C�迻�z	������"4p�� �:5x䥶MV���
2l������F�
ʞ�gE|NX�i�d�$��<.3XF[5�	�'_���ʌU����OTZ�
�ڕ#���6��o��W�,�P��#\h~/R�j*��w5~���SA�ՃL-���$X��!�H�g:�ܟ�3Y�英�>~E����8O2��^���b�錜�30ؾH�ɣQ"P{?�,������zY=3*>N�(T��-����zPRtɹ!]��V|�,��C��_�$%�}4p�{>����kS�>��̸�4j;�U�I"�s��3�[����l��6��o�U+��Bԕ�YE\=р�8,,��'�tܡ�js<&�6��-��BpS�h���[sx��P��� ���6����w���P6 �j��>����~��<7Mu����&cE� �0zf,�|'Q���O�0����K�6o*��Jb�kB�E738��dLB�aw�c����H ��˒�$�I���#/��J9��c�