XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�eLz���b�:����&,��a{r��ՁK���n�d���XU��@��>>wl�I�_���y�e�㥮�F���@N�\O�$�d1IO���MI�g2���e�w��c���_����"�#?0����"/��?��P��K���?d'�wZ�|0Υ�����^�sѺߨ���'3\OT��_I������K����'���!��O�x�`=�o*CMi�W�o>����*���e��
\g����ni^6q�7���odc9��#����-3��]�xu���q�`Ƽo�o�k/���*���qF��mG��z�t��Uo��7���V���{��a�8�d@�o��	�N�ygz�m�j�Tc��;ɡ!ko�!��h<j�
�8z>0�AP�Y�����C�φ�q0�Sz��6�/�qF���Ru�zi����JB�xT��[����.������4��B�e�	�#�Ng�i��i`)�IYʃ�ӆs���©0�t�@�	��gӃ��O�ˏ�fD��*cE�p�l!~�b��'u)n<�&�S8���0Nx���usDÿC8�hL�5���,rk}�����\5B};��D�9��a���pg5�<�W�+'�d���w˥Y��M��dᮿ��M[ ��O�aT�%��\-sR)�FU��Gǧ��*=[�lLⶰ5��K�[�)pn�d��g�ph�k��mK^I?��{�:4�g��wh:�0;[�\B�6�@|�?��C3��XlxVHYEB    e4ae    2af0��̹�8[v��R,��I���/ƈ��n��K�?�eZyt�[�f�w��8��mr���o����*
W�D y���v�aB�M(�z ��ϣ�hq�n��twy�?a���o5:�T��@EP�=���#�XE���wyGi��.h*e��#��jYɆ�!Ӡ����GZ�;�V:��� `�?诵b(�f��Ch��ZKp�~^�!�}��)z�o��En�Xi#���kvqp�/foL�ZK5=7��}4�=��� y����B^�L�-d�V�����r�����z�����y�+[|
5Ws3��l�"�f�RK�3$�.aZz����A}��{�P���p��?B��Q"��T��p��I���#�u�#7wK�Q5F�U<��<���9�����u&zz��b�M��;p��dA�Ӗ*��E�DT�B�����z��_4���<�⑩�:��)l8�J�k6�{�z���Vz���������Ȓ8�T
���#���nD� s�uD֩��d�$(�̒ݒ;dW6�����?;2��v2&�����^N]��9=c��=��^��;-rQ���I+�u+,�(Y��~�� (�m���/Ԇ��X�e���Q�Cۢ��E��t�ȩ�06�_�vs�|m~t��W�v� g	��#v6���>3��|�)�F�8h���-����:_�8�ś����^���.�]��6��0a�2�?��j�Z��Ѓm��%@�%��#�Y���~0kC�������=�er0'v��BI�_���j�iA+��!�W�S�J�.�4�]yı��������ȑ�o���*�tu[��M�"�;O.A.������WG���{���(�|Ο�Z���u���%��`�]9>�^�!�=���j������!ӝ�*Y�^M�md �$��K:&SN@�1:�B���A�s� �����ؖT��k�Zj�w�X�<$���$/��#�l��te�X�E����f�g�S�_�+]�����o1�
�.�U���\�ˌ��w�/`��{��6Z��OI��������Z��4HY;�}�,�:8��É��Q4/�����ͮj�����< mwΈ��P�����O�7#Ճ�6�>�����94����P��/#�ؒ��^�%�|��rL�\w+�dĐ����_�j��?�$8\���x�����b�?����!���Ck&�����5}�\��:�׹%�a���O-���A�Z$���.�f~�9���/����3خ�G�5-5�g�	}8 ���ͮ�Lݜ��ۅP����`��P���s�{�l\�f��_��fGO�sG�'�1����k�%K��j#˙gɛYH�Q��@,�D�nӏ�;���Z� GLX]2�7���f>7��d\R�֎LKi�����c�'z�L�]�b8��'U�ѻ����.�8�U��*���b/Hd������* `�B���pyh�w�{�͂�N �A�&�jM~�+.�.�k�_��x��*��//����ِ��C��l�hk�_�{8%e~�Z^�����l2|�F]��w��i��~�a��.g�dO�����u,E�C�:/�ƺNaP���C���e�-.���d��8NwpK!���/L�e�!l��#����U��$l/<ߑ�>H�R�_��\�CL��]Ր�`�5Δ�CaN(�o��j|� b���8ܭ�烞b���Қl���C��Rki�R��M�Ȭ��j����+�ξMMS� :=>���-R\��}�2 ^^ H��r��w�9���mk��w�@��|m��u)�!X�-��Y2.����+h~ɂ4ޝ� �L��Z�h��v3>�:k%�T�5��i������9)=\�}�p<��d�Gz0�Ìu?Ez��ݜ +|D�E�f�
'ȍa/���%��µ��f�'�[�"4�n��'�u��:��y����W��셢4	���Z+�3:����k7��7{�ts��ᛸ�7��9#��X�?����0�u�&zM���䘰��2ռ�ݓW���b� =��8�v��+{�x��E�[�Q�Lkz���i�ʄ%3�F����^X�jC�c�z��O	��rò�� ����z��eE5�Pi*ݮ��),'V�L��X"��(����V��7�^�  ;�V^����oHs��(�tl�S��
W�e���M,`ũ|��4��,|� �%������u5�>����c5lz��,j{Y��v���7�\��X�SD['�@$�lEߟ�\�g�9X��!fj�^,ɇ�h j"A��G9$,h�����UO��$L4�U9�S\�����@*�(�+��������¡	���T�̘ �v�n��GS�����q����8G���g^*2��%��e�����x�ybђU��G:p�H��m|�PG8xadnp��lJ�V�;��R9]�dʊ��
^/#Q�0��|H+��7ܔ-ޕ������ő��Ն�e�j<�"3�H�����!�$�Az�F������$$A]����g(: ܒ�K%lǤB�h�t.׾��8a�!��h��j^F����'8����~[\I��B���[�t(��o���j�˫e{�߶�Z���^W谳p#��-&����K@Q���5��L��=�z.�'	#/=�["m�;#o��h|�d(���3����@�R���ph��עk��R�\����4�cz��<qg�`J��1����
��eꛪ`�S���w��"����2�aZ��(^���Ӵ7o�F̵ݷ�a��`=?9:�2Q�T�uU�[ٛ��	b��Sjzć�d���E=�DQ��Ke���W�^/:7�N熐�Uw��<2��*�e�=�
���
���7���8���CW����RDn_P�N`,DpX�!�E[4M�N�v��B��a �X�V*��T�S�n���9m����9q4>�N�����\��D�z�ju�.|M���S[�F��#��@qo�6�f¡?�E�WP��"I�~��+��x�΋4O,�4���]V�vNh�.vvy���'�_�f%�[�PG���ڪ�L�C�D"s������ 螦S�n�V��@�1��|3��u u��bY��f.�s[8�D����7��{:-��"��(縝ϋ��?@��!p:�8y�
ȡ�ɴq�i�9�՛Oa����E��#�����"��;{�:����Iam�-#O���-�l�
zt�Z�*>�����m���3���]���7:R�^T�-��+R�5�ݏ��aC�)u��d}s����6��,�c��Fx�[^��?�e�Һ��b�M�n<.��_��y��Z@ߠ�d�s�IRg���O�sY%��;��)�܏ǩ�_���_s]_��vudAgLs���
�h)�|!����S�Ҕ����ގz�C+O	-J�ȥ8�$��X�Զ�U�3.�mWe�Q�H��d_�cZF֩"08�'Kd��d=D�ďc�@������0<���X������F�b1R.0�kB�*��]�8��PdG��,Q�t4\��N�1����=S����_��Y����p.��ΧVV��WÂ9/'�'�ˆ�xCkaԈ`n=�����i2�����4^���}b�t9���bx����I�����$���U���8��ÈL��������`����rO}Χi��ꏄ������#����f:�������S~����|[����b7:7ȧ���.���ͳfR)L��_l��U���(�����n��^1�\IP�Ӊ	IJ�='a�)qXt4KF�1�L'�n�p��d�����~^t�)�Q��<Ʈ:��|�������Y��.}�+lO��"JT�/NI���%G��_nlH�',�rԧ�Ѣ�Z��Ū���u��ua�2J���л�y&y��좇�W���w�K���%A�]j���C�C�Յ�t�mx��	@����.J�! ��ms�������?�Ky�Z9Y�Y"�.�b�Mdr!f�-i��Zbf�JQ�g_αسƳ4�8p8i� �w�A�W�
i�v����*Q�� ���|
Յ��S�7V:���i\����
襯�䣪`�&nn� �b�"�o��*����M�,�d��׳tT�����\sԝ�TvM'1K6;�5�B�{u��$����:�n �X�ԁw�%Q�|y/� �lF$ԟ��$���ͥ��&o����&�_Z/�D^LDN��ʂ:�2�'�����?����v�d�3�����GcvTm{@����r��.�3XҾp��DJ��<�~�n ��0�\��'�_����(��a��~OeKE����F5�Sy�.�Ll������5�#��e/�d�N�N�O~#�\���ÁtO_1�O`����?}'Қ0�)#peVD����c 
z`E���ZN�S��VI:<�m�V���sj|�(g�Q��T���ƟL��L1��;��x,�6�N�8�����߮>�;K#h+�)�8��I�W����~���1&�#�$�km��]����(+��</	@�U�Q�gyq����^<Z��P�~��|�[mX4]T�~�L���@�u5���e��-�A\ʯ�A,Sq=�*:�W�rGՊ(?��A��$�+�%�C� ό�m�`2���s��<�v�zmN&A�r�Yw}Ssy|�&�E��7m/�tg�/���q
��k�bG3��2Њ�^��(�.�T��6�߿��	��;�7-�V7,�\}���� A�Q�zxxf����Z3i%��$mb\\�!p���|H�K����&�C�����~�}�����h+cO��đ����j%r����7Ł=]��;�i�gn���f胢�>nA֗��<^�a��y�hdKqs�(�6`�z�x3(��o��j���p�L��q���C��=dO0�>Luˬ�H�ҙ?� ��F����2Kd�V�؄].g�D�U�����j�Y�g���=��g�@�L�
��0���˵�����Ѐ�la#D�DN}㴴�d�m��z�h;��(���U���Z3��	#��p{c#N���[O�C ��ncđt�|�̻�<G^��Dp��g�������n-Rb�jϖ��O�OVֹ�f��e��ʣ!��Yۚ�T�*�(�<�V�T���|�t�R�x&=7h&�$6�x^��0;��L��qT���F���OME6����.��<}�{0WF����sĖfm��b�Kt0���M �*��ƙ��S�N6��[�t�4���1�5������ר,����4�Ӫ	���mRh�*q�Ƴ��Cd&�P<�; �F珓�Xƚ�{`���3�Ueg?u�0eJ&̾r&;ƕ������5rX�ϰ��YѰ]ȑ{	"b�<�V���˅>7�5����N��P���#������YP�
f(GɈ:�g�����O =�[Ӄ�I��{��T�C2��L-dã�5h��5�ART����U�� �Þ��T>I��=@�B2�aK>&&��鬒�7��|:���\?�����A�,�@#��06�^��c0����9s�s\����2%�4���B�4>�X&�yB��� 5JJ�	���W؆\�,�)?,�χ\>��3+������+�B���S�N� +ҜE�{�kC"j0��Ũ�����a��ɏa��%FNQ�h�lME>`e��Pv�6��h��u���{~��DL��%�4��M8��pwL������$W2��S���6bd���mX�2/r�Ϥ`�ޔ��.~�E�RՉ�`f{���2A#���*���T`���5�5L�G�:R�9�@��;�l b����u�XN!}BQI�r�	�2e�z0�����j��m�z��E�!�rT�� gm3�ݺ��,[�΂��z���,��'�7��R6�[Q�p#���i�J]�Q�C�+��u��Z�j�:F��|��(�����"�	�?ߪ=M�9�Snm�1R�W� m���X��(�e�a�t����\���w[��Z/փ	���X�ե���N�J�h�BY[��[XW�g�H�R�N�Y�}K�-�8�&�q�Sd!7[�pSr?��ZKዥ�S+^��&-�I��tk٘��C�F畠�����L��Y~R<5��e�#���������{��V�����C-Mu����SR+�$�ʐ�zu�ݶ#�$�w"T�#�Ľ7�z�cE�z�\���Wd�G�e���ͮ�u��|�-�Z��),j�@��{�{cwjr: j���5��0/]0�8�M��M��*��E�#��BOza����"��	��)���n��U��9ԫ	��*D��1�Y���<n���i����sW��S����eZ�v��J���X`nSP���^@��r�Q��m!����{����]�U�Ț3-LM�
�"�a��B�z��aخ��݊�ǕacxI'걽dA��H��I��b�����9�,��\�0[x;�ZS�5h%$3��0'�/�^g3Ш��q��T{!XRM?�%��{�K�rX�o_qڸ�����u�Ʌף���2=u����唍��c^.B��#:�޲r.#��b/��`����R��=7%C^�N�g�m�w�@Σo�,��m�ȇ{r:�ػ�>?�ˈ1H�w��{�l��&��� �}��Ż�
AKp�\#��凋�DlS��H���J�}����̏�
��q�+t�>��u�/ռ�`)z������f����(�$p{���m�� H�_���;�/�y��˺A����� �M�w�1Q����UA�%#+	���	���	< �Y3+�j?@����e�X�n7���1b�'�1U����E2�*���FЏ�:�`��uz��A���*v�ULm�I���@H/9[�w脳7����-�܏y�%�M���JK��e�;Q���[�2�f� ����R������c��p�V���-��$�6t���m���k�k���*zEP�����s@��n�� �t�E��.��OLmK2��cPڜ��w������b,�"��)렀��^��V;EJ ������.aM��sTRAv SM�H���8�K����~��-k���bw�)�vL����K����Ds]�QL��d@�"P�X��i��`c���\j�ī���}8T���'RE�(@�2]���vj�ʛ���*y'��p� nUա���w�����ů'ĵ�2(��+M��:W#YJ�z�m�`�;��t/m���.�gM>�7���9��N�=C+�Sޖs��f�Y[Д��TT3�ف9ֳ=G���"C�CA�*�:�Mwi�'C����z��0���|Rͨ�Z]�6�Dtn���l�yA�&u3���[���j���W��w�P��#�nH=���dKu5wl�2b����B"������>�,�s<�pذ��N�g.<�#����
9/�th#�߈�h�;4���1JJ�̃�FZ��'h��t��g��(�X{m���[�w�m��-mU����΂lM��NS�O�0.=�����tL},�ռ���1�;�^��|�͛e��O�g�s9����c��4��M��V��jQE�a�t��[b���}F�Y�/pB��캆AË<0�c+$Rl[Jn;�I��d��c��	������=�����զ���>�L"φ�k,��u؆��
�3�I���+01�L�P�\��,��$f��~*��;�i�Tm�Lb/�t�ŀx�g�vC_v��J����]��⴦m[��l�	��\w��zC@���2b4���:��C��J�}��v�j�w��g��!�A������ڤP����xc�̂i_9����"���!��K�mVHn�������_:���!�o�P��|%N��f,������SM"k\�:<G��f$�&�_�3d��8k��G����ἃ����^�Q������w<y���Ϗi�.^��z�(��K��}�̹J�|%������"~���$�!�������Q����ϒ/-ϨP�|��Q+[G�1l�� �C����[	Zj9�m�R[��I���yT�6�ic^q��V}����g���b�I�W)]�*(���"9�4�L�u� ��Szϳ����C�Q('�T�eDL;X�-�hv�ѣG=��gu��_��4$�V�����MNk��I�tTw�5X���%�.n��LMi;�P�8��!��j�t0:��͘Ǌ�����X��]�=�o����ʣT���k����5�����(іB_��k�!*��쵋����~�"��4�=o ���T!�C�(�����%z@&��O\P�E;�f�%�����)�U�T'
���,�VU�)b���R����Yv��K<���!����˚ѣ{�� ��73�!�9�b�tu ��1�bLSI�`K \�������ݟt�u�(z!?HI#o��g��ڎٰs�nȃTbg��g��8R�s<��n�<�"�B��}�Xn,M���j��3��*s�O�2C��oX&�A������!F_��e��ͿR&����b=����E��t,7�:�@g_��v�E_H��}����b��Q����a^��޴Lx�q� ���g�L��/��Tஏ���	E"�#��d��T��>�p�'r `9ek�1q�8%�Ov�N�\��٭�vg�ԸL��X���¡��Jì�e�}�c�К���\M��'>ԝ�6
<1���K +�x�X���K�;�,0u�=@R�� �U��"H-:���R�8�	
�ԁ`F������E�:�h,�S]۬%���==gĖ>���Kň����|���W�f��]��\k�%�ѫ١{�}L�L�l�O-�]�N��wR#�d�)(� ��<��x{�<��%��	�MP	��kc��$�ZUT����-N�����ұ�����x�1MmN&�]x{=��b	��uՖM�!���M��������b't���i����G���dj�Oo3�g��52���-�Ѝ�Lި������)D��߆B �cq]���kؚ����c	���K$k�x0�fɅE*4��˛u�/T��0�
�c�6c�]ǜvUc���k6��� ?��ڼ��#&$�}�ׅ:�7j3k�ӺC������%Į�}��6J��
_���e᪑U���d�m�GCf��Ϣ�4��$�V[�S�-�w�����H�P��]A�����D����t����1s%�ʃ�˂V�?�j�iqfU�{�r��<�{K01�
�R���c�M��i�:֏|�<�b��#ZX9jk���-���R�������z�`<U��o�$Hz�����+�N]BAN��o����ȫ~l�/n!1�B��3̂Z\4�)�� lw�VU��8��)];�+��QUT�WI�얾�����M ��~-x݊ޏ6��}V�[>��^\��7:B�s�)( ��_E�Q��AJ��U��\�\��}h�z�T,�������Ci��6OD���L�x�"���>�����lH�o��,��zS���)��}��l�S�֖-�N�Ǣ!��_�y����ą�������0
C��N6u�n����G�V_|�w�L�����p-�ԔPU��t0`2���+a����à�0/N�)IR/|��+� f�~))I=��_C��E�r	J� �!]����7���R7���V��l�{:�h%_�{���E�jg�=�|7@r ��i�u*�/=��T�:�z-3P�gy����-������|	�Yv��	�L��t�$�!H_/�h6�8��$A�~q�J���u}ӡ��At*[� x���a@�cFA6]�iO�)fi��"%Ͳ�eU}�j���_�5�U^��g��6���\�.�d/�{�ۯ�\��(5�F
����o���C!7R��/T��ȴί]�*�#�=2����[!Z" �v�޽���TQ~�g3����A1�c��:�����e:��;���̙�x[���g$�;���,T�ڑ2��(��"đ��#�cq�W�˴��Z�/�,c@FvL_0ݎ���.�����t��z�E��f�ŉ�#D\����0[C�����Ӌ�C��r �����O4��yl�E�Hz3�[��ڋ�t93rC�6�_a>1�!7C�S��+vۊ�x�������l�S�8�W` -!�Ϭ#>��~}^��ˁ��q�#����?�(K�,�����=��V��6���En�-��l���M2��CjA�pcA	d�*�!175���Hl��$h��n��iCUk��Q�L�T��=�/��Ė5�YT�e��Ǫ\��ڂ��$�����JsDm�����w��ڂ۠��f�^{$ݥ�ȝZ���<	�����G�եg�yk��,
���_��=��Ι����/�f�!^��x����J�P��P�p?؄XoTb��^�d�0��Ma`X��N��\�3I��nP6��˛�)�QFc�Q�Z�V��GE3"۵VR��N�I��m�qB��k����@�k�|��>~
<��	q�q��"P�Q&�TNխ���� 8^G��T?��pgW�IW���H,\�a��d�a������t�s�,(B[f�q��H��d�8�"���%�����xE@��a�f�\�U�VE"�9�N4��	�h�q�}�Ib���vƝ��|��|��g�c']���4Owp�+��[䡎o|0����LVd����j��h/#�� r�|�Ŕ�
���8~u%H�,k]�UJ�\��HI�9ı`�y����o��-�݊�'�Hv��q�y�S�a)���4_���j/x��2U��MǄ��{�ՇX3�2j�P�<�5<
aRN3kC