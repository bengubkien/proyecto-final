XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1�P;���{�F^ ��X�,�|�1���3w�5�^<�vŊ�F.G�>�	�5*�R�zq!,�ډ�(U��f��>bH�^6T��z�dۂ�Y�N7���|�=��1�9�L�����[BW�?�{�5��c<���W�F7�헑O����0�l��"F�	Q�6usj]�6d����LJ��&b�S�3�܏�k9y���vچ�3,�\��n�k��Ej���e���9�t�`D��o��Ջ&TGh��}ƛ�ˮ�P�:�zb�`��C|���Hd��hI�:�{YC^*w�͊��ayL�Sd�؍�:`+ �Q�aǠ�\�v*����S�j�|�[T�eM����4�\��uf��y�`���N�':�^����M=l₻)��%k�`�H(�5x�eFCɇ�Ih �d��&����H�C/��ǻ'�+q��6�6�*�Y��",y�&GD�m��*~a�p������E�)i"J��M��-@UNU���1��T��<���id¨��*�p5����]+w1�9�r�2�e��iZe�l�1����'��QuĔ���m�S8��4F��F\���)3��|�pe��7�l�0�ށf���}�[jD�a���Uo.��3��R9A2�P�=���a;ihl�f��(�@$������ÚvT�Y�ԑ$e�"�+�&���B�/�]��L�L��[@|�9�����v�b_r�RD��b4 ܊�֠>f����]�e�"R�JM�ȭ)zXlxVHYEB    8864    1770p�L7�S�S��hO �J,Z�,���iR���s��![ѻ:'���o�}QO�,�M�֘��F$)pU����j�6UzvO>���5D�F[��0U���w��ҿq�63ڭfy7����q�z	m^̎��\�V��ث�����B�[��mDjQ~EF� �Z䨏����q�L(]H���`����ěl	��d��	�c���U��t��~ѯL>o/�s�j�mS̭S��_��?���3��'�-�ù!��P�ۊ~f�Z��+"6�q�WG��L��d׺ҜO�y�ťo ^�؆�2�3��5�	2T�Lp�u�XÂ6:p5jr�@�� �\N��M.����A{�W�u��k�;P����fx07����KJ�����`��ţ���j��!���8ߨN&�]���7?\�rK�75}�����_��x*��+�u09��q	�!�6+=T�%+#�d�/@�4�y��`��g����;�d������v��#�+s�ǌ-҆�ާ<v��=�����]70l��.>$�����4�2�3�/�ܜ��Qۘ�{ZY:�u�U���/m�- <0������6d�Psv�����_ɴDX�v[�=Tևk�j���6u�S�R3z�<|j���u�l~���pQ#�������_߮�25�"Q{���1aQ�H�~W&T��!D�*��ތ#���x���Ҹ��D\��a2�%*��yA[�@a��J{GSo%�ݔ��DԩLiHQ o��:a��w�2�Ђa��l8�q�ʦ6�ZgPfK�Η4��r>A<��<�X#�^h�m�j����%���M��+_���qٚs�|Lp� �$;
�cÿq�?""�3��e��{��'��ݫ��}���_���x�@n=+���v��RI�`���&�6�� +���YAEر�+Sg3���ЖU
����IM�Г�N�7�A��n�զ��-�o��S�r�	M��Nz@3G�w�Y{y�����5����sP��$��J=�v�Q۴���a�5m�y��V#�N�(���p���^t�P����Y'ap
��&�<B�$M�Ӎqkb���ɴzZ� N/ћ��opȁ��J�Ʊ��:����rb��Xm���u햠dH����/�O$���!���P�^�u���v��r�+I^�^0,���&��sX�.�'�� F��SN��ܤ�"��jQ�ހ1mϽ�V��s�� �^����)t��G�GjPP�r�����)<�93��Л'X��l	ռ�}���w^T��Y>�I�W`D2��E|�h��<�?�rch��^�E["�_#�4m�jG�~v�f���F@�Z�Ѫ�(����&��]���D�ȩp���-�b�#�a�{�٩��?/Fռ|�6���hj�(|c�;G!�Bayo4�>dTeø��aB��-~C� e1�0��}m!i~�[g���(�8OR"����Ԣ�I���ݝSr�;�6�a�����d�wGBA�/�7tξ׏�Y�q��� k"�1��W��"\�#�|�0+��dɂ��P� H��3�)���ġ0{:J�"G��ا���d4� 3=�#��9fJ� �e;�O~��6Q`o8w��cv�]���/FG���r m t &4�o�Ʊ���#�sÞglf�#���0u���@C;�]�"���t�v{�}���!��g3�bGj�%6@��5=S�^Cw3�E����DE�M�Y����W��bg2b1#�U��0���6��Y��^Y�2��X5�kӳ{?Egc��j� ���3�4�rgT�,��MS��G	 |�K����Ϟ~י}-�r�l��h� T��_���m�(��NZV�*��2��5;^N�z�a05�-���u��k��� �ܤ�ĄS+<K�a�:D��q'#F��έ$.(�	�߈j��a����<9y�DK�����6�D���g<m�շ��ǘ(�cTi��h����Icx��XS��p �$�������n3{U��W�-e�t��TA�H���}�zR�߳m�TcYT^W.�t��A���Lts����+2,A�a�6n���bJhN-~� �:G���˳������T��-�5+��_g%���{�-y�Ԋ������x���Bd��W�Fd�
�{�l<���|����:�����O��';�/�|�ON R�YC(ƃ���k���y b�ޝ������.�>h~��F�j�X3��\,�"��#����/1���qIWͅ~!�� ���5���	�0Q�(aɅ��^���?��,�q��ɏ�R�"J���&�\>�GP�λ)�G�l���#U(E�Z��d�ǿ�=�)t��H�x�|��FrYʡX/$��F�������f�
5�w�u�*x�9�H����y'��f��4ߕ�x@Q�-�ge�*K-���Xpq_5�59E{�E�3,ꊐ
�2*�	�r6-��M��hXO
#Ȑ�g�����G��	�/�������a�: ����v K�t�����$'Qe�q(�h o*��n�D��q��x�^$n�T�|:w(��v4�f�{�T�Μ8ё@���*GQ��Rۚ�xW�nb�; E� z��A;��y��B���F����K��@����Z�D꫊�����64��_S�9��s��9����3N7�	oΣ�@�7V%��잩,��bSC��͒�R��(�g �"Y~o�\�id�>�(���v�=^��ǳ�۬+7d�P�H���g@�������[*�M�|���X����!yIV��$Z�]��3��8�FҢ�!$��j��1��[��htH���	c�$���D�U	3Y��=
J�ԫ̤J-7܌؞�<������RMg��׮$�)�� ����::������w���k��J�:W���i� t&$�g��_ƭ��?�f�1gq��L�����0f�	�O���7�@PZ2�K�o��ׇ�νi��ʲ��/t��A{'�J�C�����V���˒Jާ���G��!z��il�2P�4�㿳EJ]<�$�
�".��OX���&f�x�
�vx�3�"���ƹ��Ӵa��[
��*'K�f��->fȎ%>c7�� F�����4eWj��w��7=A��|Jb�!p��>,vlR������@��DY�CMC��ÖV_���s=��w�Ճ�}Y!@��M�7�o:��Q�)w���QY/�cP�fNE��P:�F�/
}�^㸞�MkG�|q8�1m�達�-�W��K��'��J�cW����<ߏ�����qa�{�T፥�xiĞ�������朋$��/�X���k�k��	nX��l,���
�j����^J�4���=���UL���K�R�p�
*��0R!3�R�T�c|B��g�;<$@��4��H �)�-�b��IݖSuTo�[Z�z9�F�>9CK�6�l�hmdp��R?֌0~�Yǎ��X���6�ii�Yv�X�q)@�`�-uG�\S�d%�6v������BZ�Ϙ�BDYA�I._
�7H=�8�������gy�zւ�2<=%|c�����r�P;|��qթ!��̤���'�`��%^���_F�!;���f��*(�&1�x�=W��2�K����dB�Z����1<~�R�i���s�C���N��Q��u {bqB�	��:� �[�����ލ�7}�MMCZ 9��_l�SK�F��_�޹��ęl�/�;��%6���Y+Rd`�r�a7P�����x�.r�u�YoB-��5W
2����7j,O>�ԴQ�C6��V��0M��4�8�(�`7u<�"���״�Qk��c�(��A/}�(V�`���AR�E̸
h����8�b`��Fy���N��B�E2�A�~�nb��k�0J:����zWMG��i
/gGS���D� �j
P��]�ݹ#k�/�>X��lPg��_~�m�K6rB�����ޘN5Aٜ����;����85�:W]�ڥ05 �� 2�%d-N	|��V�[�+���`w����Lp0Zܾ�U.I��7��"Owx�c��o��{�T)J~�l����Q!�K1ׄ���-���Fb�qv6�4Zlު�݁��)Q�#�w��ܾ9�,�7Yl��\���X՟�fԦ;.\��,G�?Qy�`��7$<Q��֚� ��H��cJ�U�eK��]4B�n ��!�&���v=����uŭ.]'�Q���i���.774X����D���PA�m�g�l"l�,:MJ>e�]�h����Y1�Nq�X[���vĂJ��!�	��z��{-0�خ� ֊_>C��͸�_;���<���� �qP��2u�~���R$l��B���Wڒol�ZE	�3��
����^��3�0�A�|��]d�~�:5+�C\e�/T��FĀ���.=#�<Xl�!l�H˽!�&�v�"<��:A��;"xe����� �_g�}�{l����^�K���K�H�@�����<�Pӽa���|���~���}�$���ɰ齭�%d�c�1���U��N���W���Jg/<<�� L�Y8y���CR�t���N�50c�,{��1�闒�U��T��C��X;j��c#�F!�{+s��Vr7
��5�#�j�j˽8��}�_ bǞا�s�GN^����f�j�MLr'�)<���AGY�Բ�9:~�"�f�z�̥]����~��4e\�C��w�B{n����/٬���$v�'巧N�aE��n 3@mCԺ���\)sx�9�N�rɆ\]d7����9H�A�������p�6Ů�h_r�?cf�s;D�T$]5C�?XC��ԟ���!�`�^�I��֟8�׃r�f�?L��v(*tɶֈ��"
#Eeۦ�Lh�\�~45� ~W�b��!A�$+��*�	~ ��q��_� ����xi�=�t��E8��^,mZ��[�O����)����Ru��$^��!�-RȪm��z'��mŧ�E��D�����@�"Mj=�	��m4ծK�2�Iॳ����["�,μ�Af<	�F_�O�Q��# ���Ѹ�k)1GJ��w
�8 �ǎ�i'���z׎�9CI�BjM4�Y��ޓT���Q�c�C�����7L�;�]JG�4��a+PS��oA�ڱ�����ؔ��3G�eD�r[���yLV�T��G)�sk�1zO �?�o�Z-��l��Nｍ�H��bĉR�Ar�M�'�������`��6�/ ��O��B��8�H�����������P���r?�EH�T���:<V�t"<�r߫I������* V�)����zd��J|�J��W:X�j}��+�i��3K)Ŗm;�Q��?�����TV> ��@�d:E���؅||��1a.�H�WL�%:0ęe���I#m�"=��]x9�e���Ya	���M�՘�圽����pD"1OK�d�˝#"����&�w� /c�����������i?�2�#��n���!>��������^T.�$�d�*�᝼؃�$�(�%?�����YN_��:@<Y"8$�"�^��_��f��~��^�6��8�4=y��+��4��j�~얪g�E-��8��kH���>x���6����Ю>R�Q�q	uQ^�#[F��>p��e���gfv���w��|[���u�oL�0���|F�;GҘ����0�/��t�DH0_ fӟ!=�0��jY�I�s�g�{��{�m���[$(q+Aj���ȕ �`�$�0���L������E�fu&�������#*�_��״MJ�<&�Y����߉�b4������=��/����Y|�Pz�Y��`7��l�{��%�|ו_.��5�ʊ����Z���4i�f��K��V�๾d#�;�FL���Q����������f�(�+�������3YP��;k�;��ݠ�p�mV=CI��
�4|WߝV~�Q�� g�' �����xe���\^�Kg�=Û�>�*���	����Ӡ�k�9���Ä[gL�