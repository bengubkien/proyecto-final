XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��TW����W-��B��-�`Ǯ&c&$y�������P�4�c�ʹ�UԊPh���AW�?�J0R�d�-�8˺����np;���]��U�x ���s��=�����|\V��vj�;x�M�)�L$�i&m�x%t�.����״���m?F�08R�ej+(��K� ��I/��mb�+e��5�O�DO�$�+Ac�&P�
�r��/��>`Mʶ��.p'?6����ta��i��x=�vˍ��"cO�Bt\奌��=P��VLȷ<+���Xus,D���fW1j�"t��6d� E{����b�2��=�7ʊ���Su�4p��%Aj�a��x�hJ�)��xX�M^nfʻv�x9��c�w{x1�8���m�ǭ4l�N�oW�������Q��m�H�P	�/ˀ�/���X���*�9�r=O��9V�씝�_����o<���׽�5��ɒ��8�E�W&dl/�-e__�(�y+�sD#T��p�@��� dԕhbЇ=���m)k+�g���|��%�1f�H3S�X�Z�XZ�	��G\�7�f&qOyhoЄ�J͎ΠJm���`�B��j�jX��1瘑�	��(Y�������H�qB��^�1<5����<7�5��oOT��Ś(���۷2�r�l�1����%P��& ��B�3^�Ј�Δo[��6����.�T[�BS�j�d��ts��E蹄blS�9�Iv�wJ�Uy�G��J�e%���Y#��f�j�j 7`;	�1�r7ң�<L��1sXlxVHYEB    ce38    2800i�dU9c,�Kg�yJ����&��&��O�tF�R_�a<�~w����t����H-}�Cپ��ߎPد�K ��.��`�g���s�(�R��çߚ�d�b�n�q�v"��le�b�hGL��݂�D8��2)�Pfz����1b/���3U���\�$U;��1��MѠ�8�e����Xc.����k�ő�	�	#����Y���Yk���c�_���w�2H�Y&���W1_K�9:�`f4��Q�?֫^�'��3�L����ն�Y=n�0I8����e�86�}>�&�N��N����~� e+
�DR�\�%0��P=�hI�z�8��-�A~i��^\�G���3��!����-8f�{q���S`f�N��Q�qͿ���K�
R�+`�M���M�{sܾ�?��ϓQ��F֟��4�]}p�-�Pr�7��A�M|9h�P7u���`�s$W
BG�R��UE��[6�z��((`��S"5���/ȓ8���)�H�˗|�.y���f<!�I,��&��`Kw�N����>R�8?h�;4��)���̙�6`
dd6_xT9wi� ���W�)�R�Ql.	z귕�>��mk�}��6nX��K�+�����'_ąLVe@���?Y�>M��2����{p�=6�qCD��Lvl�n!�M#I�t�I$�2`M*�U��yF�$�9~
�>�h��K�X�5��4�C`�5u�Q�2W�zp�]^��I��9]���o��)SH���[�l ���GJ/����n�P�؃/uGlj�Yc-�b�Q&D�)�pn��|�MT	��DAf-'@V_����Ո��1L/�` ѕ!��~Jt���?������s��=�co���W�z�ٜ0K¶H"��K���	<��a�|���e�2��&\��J
�pxA*iZ���ڭ!E$0S��j]�M������ЮgK�i}�}pѤ&��_s��0`kA(o�vh����Rs�����I�����<�3JtY���T���2��<C�KU�e ��0����@@�S�dxV�K���z>k<���&绝��P�|�Z� ��ʛ��4[�,�ӟN��yKs�g��3ӕi�(�v��^Ցlt�������}-�y�Uѽ���[{l����	���|���H8�p���!��|�,��:�ڂ.˩I4 �X�y�<
�Ι�7Zvx��4T.��Q�2�4?;�(�� V���M���F��jSj�%�N�@���
%̹εu���\��7�%HL�S�0:���9zHc��ǿ&	��f�$������3�������{�"��CH�d7%x/��o�ݘ��G�B��,_&�OB9BM�_y�.l�Ҙct��d+�ùN��OvE����+ԀW��M!�S�,�
6%Ot���l��lt�C������_l��t8�W,��b�T��d26f4�޻7��bYB?�v���W�3��.'J ��1�S��I���1)�w�h��mI6�i�k�t_Y赣�`��D�4:��"8������%�R�Z7O?��s˕'�V��>�w�J��N8�n+(���=�q�i̚�c����3-��B���hX�㺪�K���:.���^��g�v@��Ab��{q����ZR�Bo�1͞�Lm����|]�;�����^emE�������wDƷ#fQ�I������b�8�Z�#[��mK�E�vǚE�P#�ͽvP�K'�*2�64|���%����{䗗Äƭ���T%YAQ�r|_
�Fx��"~W���9e9~��*��tY�3����"��{�Q\`�ׅ$�U]��H��D�7d�I��}&��c��C%���P)�����r�+�n�T�2O���W.��6y�O~ml�鱥*��O�(�	-W��o��y���@9K��prd'"�"�G�,b�=���8�Ά���Z���Z�'�� �c���ַN�B�v`�<L�G���Td�ɰ�Zf�4,�������̥��kcq�2G��x��֪h,��)�i��J��=ͨ���WڶV�e�ͅ��H��,{�R�;^_�u�]����+۞���ȯFs��Ӿ5c�RP������k���}Pu��5PǾ�x*���M<�Y�n������V�'-ۜV)}A��?���<(��*��=�-]�.g�&r�n���':�ܷe��ZkS��yS���.������G�ÉY(Y:!�%���#�\|�6�XAu|a���_��B�I�փN ���K��տ�H���iLa��M0��8W�[�7�w٩�j^GE����d!������!@�t��C�o�|�g��pq-�p����
ՙw�߁�Cb����_�J���B*��^
��egq�G�8ݔ�� �t�;��.���|�
͛Ή�d�: �{�1�&{Ш�a[E�,`�j��AӺ�C^:d��+u����X*Ut�lo���	�ahز)�8���gM��WB�O���jI����-�#�i�Cn�C`*�uñlQܣ~m>� �kVCl��Hs(�<q$��UoìCuIW|}�r�i39.�
gkt���q�+����Hqh�����f=
�'��v��Gi�8qQ�F��)Rw�`J���v~.�s��#��{Ȍ��� �f�u�KBx�����yU&�Ӵ���N)�.�|� �_�;qH�|ϥ�E7�o��*o���
�.��DE�<���	��
:��Ti3�;�ͪ�rx�G�b�J�2����_�.OmxN����J�Z��%���5�M��/��	)�*0Mrf�4�#pG�u���t��'L��1./ǳ�ۇr�{Љ<��HDAY��
�M@��ET����鼧�O�����u���Lf��j)�8�b��2��a�� ]������F�T�\qhR�W�_�tc�H�1 ��{��c���s	�� Dak�A%�+)c��I�����}��)z�V>Z =/��3��g�Ͼ#0��9���x^��MX5�`^O��uS2�r췄j�(���7d�3�Q�X����֫��%Y	.#Mn����h8���6�*�q�B��:D$Ӈ*5�E��H;�`�ZVx�M�"�0�g��g㽺�VrI������$1�.���R����$ ȕ�><u�^xs��*��E+
���hr�X%ML.s���O�<�4�wȂ�K!�����W��W�~�m�գ���7u��y�C�{Kj�	����[틊1I;�Ho{	l�DvZ�]�]�\3o���+/}F�!Q�h�L�V����T���!�v���K�߷	��6b�ț>cJ1ZS�I�؈Ct�ǎR�P2�{sǟ�=,���>��Y¥`㴑j�J������>7�7�'��X�n��}�2ɣ#1'x�1��#��"�_n]c��uIڒTe[R�P�>x�B8�Q��� ^����=�f,��m�zg������U��:;�ޗg3��Fc̊M/ �Fj�C(X�ӎ���ISn��2���s����޺6ߖ�,'�*�-���c~�D��4�l�#��L-e4K;=mvq�j5c��6�Cw�~��vL�h��Vq���#B��]�D�:lٔɾ+�8y� �ly�]��t��D���Q�7(�]I����_�/�7�7|6k�Mc'����&�2aĥ�l֞��=��)��9M�z>����M�{�ڇ��"�01��/�C�bI�p��,��S:S��VN����nb��E�^�<2������Oհ�hC�=����4<2_���t���	aC:��z�v�¹������?�좨\.��|���l.=X��k��j�
��ң��e�A��l1அ�N��atF �<�_�q�ݿ`��w��]bd����$�}D�m ����
q=��ҍ$?��_�d-�i4��@ԍ��	�ن"��:V���d�R����N7�C�0�Q �f��)�mQn��!= �w@�=�e|!4{~7ɍPɓ+���s�*v0U������-�}tP��ڹG�я1uE�ޝKM�|#ց>&�f2^A��㉿	pо�^Ju��]��8��8�X���d��{Ǳ�����/��/��M
n��|��-�*��f&���m���	F�C�]M{�?���^O��a!Ĕ��2�lЁqw"(C��:8w��)y�]Ҫ�[��;ꑗ�4)��lZ��O��HWW�Z���{X!�������ך�m�.��HX��t���PH����^Q�4
��Ɠ����$�o sgD8��5���%$���>���*�Eu���x�^ہk!
�'�v�h�)��h�+٢����0��r�p?�s3�^)�������|��i�B�]�X�e�R5tfE^h|PKP*��H�,cj)_$i�LTX��OiS~����\{�����<ڗ�w�B�pC�)"���/@ό�rTdC���wDj��V�e����)7Df�;�2 �\�#���,��(gǀ�̙����Y�ô�KC���Q���������ۄ�eՙ*Bke�*��k���wv��8v#��fp��㈼���|ɭ5�������5�<8�����Y�n�4��^ �,%�F��f�hHBG3ۮo�b<O:ޒ�|�*KH��f�T	C��\0���|=1�C`��(�����ca�w�ڦ�|������Ǚ�>�-؋�,O.���'�^�=}\��J����O���eu�>����"���������qV��m��O^(�	�ȧٷ8u3W�r����4i��.�$.�;ȟ�!��_�H� e�K���D|=������>��;�=y��lR��tX�Q�}�g\���J{�Oޯ���T5��ۀ6�p̯�־Q��`6g�:��L�E�v��ͫ���0����q��H�$T��I��o�B9�B>Ъ�9���v8l�v�-�!VA�'���� B��Yz�I�o���!ޡ>�����,>�v����V���se�����277���|Ť���*�&ĝ��#i�q��d�D"�;���͞+�ħ8
"�8�]��/z�g�I$K�.��Y�����ES0b�^�k��;�U��)d0�t�Sg[�HDi_�;Lկ/Z)9�a沚d����s%7�
�F����^����y<^K_�&Bvd'}���waF���{u�n���� �s�90 Ⱓ (�:���G��p�B�S\�e_����q ���?FD'W�p<]YR�}a��s:W�+��]�PH� "��81%�ʾ�P��o��TK��p����S�KoO���u�����$ɬi��)%&��S>���v{����N����������!	,�J��.��l]�i����"�o�z���'�A�HM��Ry��~�W^]���}���w���$�:
�|	+���ۙ��u4��m����X�#��H���]_��q��/zY�:�(�.�b�m���?&Q��8j?���C�Kz'��g�f
"orC`/�=AF�0�u�f f%��IA�m����z����� *��.��;��n9���i 87Ct�
=���l�cs���e���+s�eQS���L��+ㆮ������O�M>�ތ�����E�K�O�S���t!�	v��?��#���Vu�w�����(����Fʦ~�<��S�_2S���h�>�ّ�\H�y���ػGl�u���q���@#_B&���N�N߀,f܊�ȕͼ&c�t���tƚ�4�,P��,����W(�C�ҍ,�`3��Zp���b��*{0wa����7zjp�^_Q86''�*K^U���@�x��؆��mm㐡}����}��T�~n�i�68Ʒ�k���|0I2���3�T�¸^6�&�ͷ�&m�4�	'���Ա��W���bh�'�mߵ�̴��
��sm4��`H�\%�6�A�j�&�ʸ|j���t2�2hK"%�+Ȗ�\!{*o$<z�m?��k�S?�^��57U�����C�@]��c��U�VC�,q+����������9�V�S��m	j�����^�����a~<�P8|e��9˨��G���S.�	}�y����)L�@اŭ�_�HϽ�9=K=�;��e�J�a[����%�=这��`�w���Y$�,P/(�C_�K��푇�Sb�p�9%��s�!�u|1.�G0L��r�$r��eB�AF�B�ϋ�&Hm,���ݸ�	�78��z�^A{7��|W�6�.Z�2p���P�N��^����7ٴ��IK^��������a�t��¤ 5����I���l(��y��G���{�PS���>�;,9vajq8��a
�Ej�&O�6o�	�T��8�줊����#|�rF��kl�Y��.�HJ����U]��;���,��&
�9�2�	��}�\������/�w=�|�!�N��L�ǂ��hn�Bb���{>��FL=��-����6������nU�!��/;C�+8HIG���o��Z��FTPM��!�h����f%�	��.�I)���ڵ�W_ �2p����ҷx�-tH"���d�V��(�[��$�i4�F�Y�T�����4�-Wf��U�2��R�vo �xZ�K�%��9������b��x&�{��>�P85c�K=�,4�R8x���W���,B~��L�������Z	B��Č�M��=#[���-��C�
�:�:q�[Ts 6�j\�a���`�+q1�.��q�4w�RJM6���[����dN��&UБuG�]V���c:�M�kv�$x�B8O�ؠR�*�p�o<լە��n	�<���-8p�%R9y��o�j��#�������R�P�5�^�^YAu����
�ا3VDjL����s�H?B��l��5k�����%��*�x�x�#ȍ�O�-,����  ��U/TL�����p��<b�S���}��u�qb��Ԗ�6���0����7�>�ݭ��8�N��<&΋>d<o�\�|�b�K=(yQ��W)vY��O/1����`J|��X<�+�`���I]��V �H��l�;v
��U�>�2|~�(B ���fG���?���?�n  8�����BT� �"���^#�h�f�x>�������P�#J��1̹h� Ck��]�6  9X��c.�7�w[�< ��!�{8�B[�~��p�śI�U�j��z�M���kĥ�]���M�Ѕ��� K��� {6_�+t�3��6�,3W�i��>�!��Vz����mi2��w��7[顬��%v����=�_�x�R�6�}y�~�=s`:������*J�~7�XA�KM���"���3���C��m���VK������|R�@i���~
(D�o@D�S�ic���qv�X�6:c��ŝ ��fT`�z��1����[�� ��x�p�@R�Y����P�'�g�Xu!"Q���9
��$0�u.v{�I��ݶ� e�d�fد��K?���{������Xa�xb��A�lJ���Y�+Ryn��B-V��o���ˌͭ���uC�@��kŖ��0�v��*��i���sm��(�a�+
���h����H8�~ї��Bf.��4����e�������}p��)�Y;Q�m62t��DV�X7�����{�w���������tO�s�g"8YmS̿��mS3��A���>�vhz`%A ?E��M5.����B?w�ЗH����4�HQ5^;`���7��A�#���& #օڦ�̓[��x�MIN��;JP��<~�3Ko�������6*�h1''g%/�l���1gy�T���Pv������AT��j��׍r �G�]8c~4�I{[�s4b��+�ιV�v��	� �l4�oe�[��SS�yܐ cN��Np2����6A.[$�Ifs p�g��ʩG)~K���T�>ܸ��._q�c�8�k��3 C6�6S|e�P�a_m�.3%Mҳe]�hc��-;LV��&��w�����_͝40V��\d0RK�b]ҁڅI�ͻ<MQb�^��C�M�<���ȁ@�a�0i��4@y	�o'��>�A�ڸ��u�G��@�G&Z{��['�w������tH�X��D�Z^��0�|.����;��ޚC��p�O[U0�]⸊.�[�iSx���b��C
�t�_
T�qM`�L��S�zI"*�;G�HZ��d�ݢ�_������p�=�*����$�˘L����p� �� �?[m��(x&]`��2�f���[�q*hq��B�[PĂ*BL�?�9�P�����m3��Y9~N�~��XqĞj,�xXط7S �J0\	Bo0�2��I6ԚŸ�C�2b�l�T|t7i�N�X�����B���E�Q&�I��"��G^�N���[P�����&��:5�W1kR� ���Q.��d�se�.�kY`�2��U%��ғj�t���j��8c�Ǎ©U�}%0EY�3B^���b���@H�4;�[�d�{�*/B��@D�#c��o�p�L�\'lA�x�h@ɺq�L���*V��
�_�|�a����]ֵVi�^T��X�x7匀Cn�xM�Uo���kQ?Y`��4�N!�Lj�*>�z�=`�>� ��M��g����/��(�w��3R���DrW�\����X�Z��m�b7iX�d�Q���x��� vCh.�h�������e�������������|a+{;_Jx���ͪ�@��5�ܛ��N�b�m�&�p:��p�n��;K��TaH�!��@煖{}�4q�x};���'h9�M�2>���k!xB(}˳i�n{K�zD�����\��E&z�ܤ`��� ���:���Yi�76�"��<Gq�w{G:���R��TD��.Ѫ�!Ѵ�L�"} s!$�B��7��3�f�Kr@{���-+&�|e�
{��
|/zaEb��w]q�E����(� \6�Nւ�Q�ƕB�	�Y�x���*�9�#�:����=.�23��ނ��yI;�nZg̬JW���Us�Ә�cbT�2��@�&7Y�|�ph���j��6|�ƅ\_e���u3Si� .I]Ň�~��2|(����(��M8S5��FNfcz�:\]G"E�Y؂ߑ�	���c�x&��
�O�q� ��"
�voЬ(w��魅���]�x,���=�V��:ۇ��p����iB��3k�m��,b.��:$��j�.�f��maץ`]���#���Ϯ�������nMu9����+vGד�zKW^cA�6�k>��+����K٣1a�x���VY����:�UBn�1�m�K퓳ѷl�i
,
)��z|�e57\��7�K����E�@b^���ة��I���~g/��λ2�;��vU"��ZGQ��=B�d%�)��t�1����$��}�|��	;XZ��+C����,����t�#S!f�3��h�
����2�f��%��O�X�����ooZcdD�cK��O1|'$�sըSʐ>&�(ZO�B�4��/8���5q讁���r����s��i  �C�e/\�p�r$KM�?��>�]�s�Y�&y���ft�	��v�_�g����a.�,�l0�̆���b�Q���Y0�Ӗ��=�x��R���:��⛵�:-�"{�EW�;�=_�$�4d����V��C��E��* Z���Pտj,2��������u����Cw})Ũx�s��2nn~�b
[�w(���z;6W��o}C�=!$�T�v<;� ����K�y�%��e��]&����sV��G��Y
ظ6/UӋx!70�kO�5�@�8����q��6� �����R'/]Z0��8u]p��(�.�|�yp���;]q�9Q���ְL%!��6x<��)֯��O��:7ZI�zH��X�w�~'��q�(������5{�W�p;�m97i|����:Y��(.�S'���q��=PB�
N���-���<Y.La\�"LJs�Y�%�o2�Wױ/rqw���Rԫ�(�w����bdW�GJl�]B��vx�ԣސ�bX,��J�(���C��JJ/�n��!��7��8���+��:#��1c_�S�ya�xo���!/rK�P:]{�ʺ����h��
��-k�=��mn�2M��t��Mo�`f���2i	V���mC�N�"����ܴ�HXV������Kg��1\���dL���