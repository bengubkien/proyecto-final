XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����a/?�[+���l�v��ā;EQL��򵞒.�5� N��w�-%c�(�S�$��#s+�;ZCG��X�r�$xr\���-���E<�q={[|��įl�S%O����D{]��~�����sf8ښy ����\h�'e)��c��a�Q1�T���Vn���$R˞CcͲ�|5�����TУ���E�U@M�ф^�1ƭ��a2�9E����x�~��^9�	Y�M.C̀`�|��,�������щ����c%@xp�\w�3!���BTC?��m�XFJ��؃�h��>���d�Kd�����?���*m���8��`�L��5�2w�o�Z����Z}@���j��v�PV�^� �!Xʆ��{f$��k٠��Q�o{	����4�ι������-���ؼޒiQ>>��k>������4�1�I֟��^4�f���S��5K���ba]�H v��[��s))���ku(U��A9.�\ ��̈B���+���z���!@�MK�}X=�kd��Y;�]��,��� B;���v.r��x�U��[�h�F��B�G]�pW�ye�Bf}ݘ�.���6%+G���#��H���DE5�n:ޏ���.2���DspU���ɰ~�_�)�D���e��a�:�{fQ�;���}���`\gt?0��`kz�ue��X�C�MV����"����ay�q>{� [Wc�Ou_��U��c��>"�һ��
?��EZx��u7�.����7>�XlxVHYEB    40c3     f30ٙ�q��	�O��X^?��Z�,AJdF�c>�0��e�P�h!
����/�z�&a-����]:�A^��y������@5�T�@U�i�R���<�N�;Aߣ�4ͅ�������?�t�z�a�d{����M�K��dL����;<.�l��l�q	�+�W�p�'OI6�=�q.d�+Cf۩�po��~�d��%:О[1Z���PIu�-����a��Jxw,����Y�*�`|�Ϊ
���-���{����}u3G�ƕ�p?�����>�C����P{Ƚ>��Qb�0B"q��qEm��q3�/��S[�$@�J!�L�hkUB's�����eCM:��"���tz�5
�$ƍ7w �(�B�9:x$x��������dZ߭�*2��Q�~_�p 3��]��t�OaF�CTw������e�1�Tet���7�E�W2��Б�F�h���;�k�zC��@�0��(���dƈ٬�M�c��7�ŻT܏����9�@�5�9b�G��78��H1���K�y�<����ۓ��enrX���O=�<kj���(y��005��]�*��՜�E$G�o��.<�5�o�sp�
con�ų������w�!Nw�	�V�ou�:56���sM���@����m�,j�Nl7/��7�ٔ�z/m4_��3u� �,>R��Pr~�٣�ZZ�40�r˺/��U�/�
8=�;�Ʋ1�����f�%���fA�D)~/��"^:�8�\�M���o���#ی��,.��*,��1�+(�(,��G-�<�Vܪ
aǧl�5a}�4��X��E���ΓM�� ��1v0�Tܢ9
\���dY��k�(|C�5�8���y<�['�$��|�W�������*���x�����zcƚ�5�:vmd��aҳ��g�ݿ@?I��ٯ��Ú�ךx8����W��!��hk��.I�\+o��"	h�2]=�T
7�U`�U�>yu��ٍ jK�(�.�jN>�_I%R/pD�z��f��{cj��
^�H3�z'����zJ��\�H?F���6iY J����5 ���`�t��Qw��o����;i�쐁V�rW��/ع�5V,�]�D�
Z�ʂ+�����h���>�17i��Qp��a}�%���9��(\�B]�`{g������*���%��iR�y����i���@�A=/�oZ�̵��F0_NX��4&�C`�<c?� �"O�]��E�-����␸B���%��˛PU���*��Ҋ�R���4�6����JI+�E���z-�B(�}�;P����y�d��t%�͌g��U�í?]�[@�3�8���e�1����Y�G�+����ӥ�R{,2���K�d�k���Г�Gn@plJ�ߵFP�X�u�B<�'�5���k�����r�s9�R�ƫo�2~Q� 0|����?�-��5����2 2.�B�~�"4z���Խ!�	���:O��%�*S�
�j�䩴z��C��o�*�7�w�d�H�˛�^`��SJWrCY��*�����O��� (���M�
Dһ�;���eG9wH�����!o���0y��=�X	��1l���p7��d�G����"�����23yfS��,��0����0U7�aGg�C�T쾡�a��)1j�
��$�qu����r?���%��O�����@����G'XW�.�f����c@��~J�aŨ��"�z���f��BMl&(\098@�/2�م�*\�G+���k\�0�mG{u����Ԉ��mZ!,ؗ�HkF�?QBM�0y�2���(��7���V�������+?AK6����7a��0@+�|t`u����a5.�J�D�
�6!����[�u��j]c����|��1c��]Q��ݡ%��mJ
�d��j�I8#��l�^�3�~$�� ���r�(N���kWt"%�X��;9� p��I�5���vۨBVk8��û��N�^��^�u�dg�������1�d͊��`Х'V�s�'Bc9f*�_Q0`�lշlbK���ǕPL��u�b0�Tܢ��fU�q�Ľ
\O_��8*�r�X�� �����sX�hN����j|���1)��e����%kW{�;���pB�w!������hSӇU1�X1Xp~�u:��gF�X�?"2�`#�T4��n�y ���!iǴ���]j�����$̢)��AQ
��8���0�����L݅�0~�:��D3t@�35��6���T<?E^����D'�x�i�Z�D2x�Y�����Ʌ�9��v�鴛�_�a�u0{Iͅ3`䄒�={Y�
���o�V�s����?�a����$�l}c������!�O�̧��R���o�m�r��LW/�nG��l�7*m�1��a�0����s��i�lM�nCxc���"�	aB5���ÂD����ihk�K���'q�_vJ{Ԇ��@B�3y�+-l�"�oo(T��:�~���q6=a����J� �{D��V���ڰ� ����q�Eϑ%~���J��{oiI ��\"b�Գ���A�y����+��E�y&������P��c��<�Rp�S�o�H���
j�yP�+�;�����5��3�E�}��
sم��a��0�$�k��6H��w��.�`��"�?�o`T�[$��U9�M�{C{n�$��"�
�~<�DQ1��A�L�t�Ӧx8Xs�s���o�W���h	%����#�SA	��ɢX�����K����t֗��{������]*��S��7�	��
��F�3�Mb�
��\G��wJg{��`���ȃ����v��9�E�$���NW�����i#V�*��,=7Z��䤀$ʀ?7�� ��&�Y��,�HS�����Yp��m��������+{��w����27�x-�b�;&X2$io�ӵ��|~��.���M��NN����<�����[,nOo�Z�ܛr��nd�Ǆ��"Y�|�!�t����R���Q��I� ��m��`�i�m�.x��u�+�`Gh�z�"�Xu�	�d�UW5��������������ܾ��L�����#O!u������a�d�������-�yڝ[`U�x$[����*�!��/_W��K�웑T�T@SB�F�W,�H1BZR�{�Ix1�	J�0y.�����ښ%���#�1<at�/� �g���P��'?dKY�i�W���[�b!EH�d(�(��e���n�7b��-��ϯ�Od8�6I~ugP�eu3$t��-r�_�
W3v� �)r�*Y�{��}�<
Lh�jɮ�G@,4�:G�@�:���by�ylaԉ����[!Z9��L��Bm<k�_sq1�W�Ki�;`++o�&�F	{�y�Q�Z'T^�teL�-�~�X)����GT�ٌ�dmZ�����a)rO��0 ��c����ᨌ8�E
z\�]Mب��2�_:���!à����h᪰�MkD�6&~�i*��$!��PX����*Jf7��>d��|��2�3C���n��b��)���[[��&����Dދ�i� �*7���c.�Ќ���7���?N%����`���E.�J'g���!i94�����Q�}1S8%� [xu��6-h�w][N'����4��w���<��_�܆/t��k��b\У���y��v���T��D!G��,��n:����u�T}?�~(pTW~��K�lNn��:y?���(��I����F��_S[܇5C�*�5Re���!=�s�p|��a ԫ���b�P����i��];�筭u�x�Ŵ�EU���;f-ӴĔ|����